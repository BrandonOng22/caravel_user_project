VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO flash_array_8x8
  CLASS BLOCK ;
  FOREIGN flash_array_8x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.275 BY 25.530 ;
  PIN PSUB
    ANTENNADIFFAREA 8.916200 ;
    PORT
      LAYER pwell ;
        RECT 1.430 -1.860 9.360 -1.430 ;
        RECT 1.430 -9.110 2.110 -1.860 ;
        RECT 2.535 -2.830 3.935 -1.860 ;
        RECT 3.975 -2.830 5.375 -1.860 ;
        RECT 5.415 -2.830 6.815 -1.860 ;
        RECT 6.855 -2.830 8.255 -1.860 ;
        RECT 2.520 -4.810 3.950 -2.830 ;
        RECT 3.960 -4.810 5.390 -2.830 ;
        RECT 5.400 -4.810 6.830 -2.830 ;
        RECT 6.840 -4.810 8.270 -2.830 ;
        RECT 2.535 -6.160 3.935 -4.810 ;
        RECT 3.975 -6.160 5.375 -4.810 ;
        RECT 5.415 -6.160 6.815 -4.810 ;
        RECT 6.855 -6.160 8.255 -4.810 ;
        RECT 2.520 -8.140 3.950 -6.160 ;
        RECT 3.960 -8.140 5.390 -6.160 ;
        RECT 5.400 -8.140 6.830 -6.160 ;
        RECT 6.840 -8.140 8.270 -6.160 ;
        RECT 2.535 -9.110 3.935 -8.140 ;
        RECT 3.975 -9.110 5.375 -8.140 ;
        RECT 5.415 -9.110 6.815 -8.140 ;
        RECT 6.855 -9.110 8.255 -8.140 ;
        RECT 8.680 -9.110 9.360 -1.860 ;
        RECT 1.430 -9.540 9.360 -9.110 ;
      LAYER li1 ;
        RECT 1.680 -1.730 1.850 -1.560 ;
        RECT 2.075 -1.730 2.245 -1.560 ;
        RECT 2.790 -1.730 2.960 -1.560 ;
        RECT 3.150 -1.730 3.320 -1.560 ;
        RECT 3.510 -1.730 3.680 -1.560 ;
        RECT 4.230 -1.730 4.400 -1.560 ;
        RECT 4.590 -1.730 4.760 -1.560 ;
        RECT 4.950 -1.730 5.120 -1.560 ;
        RECT 5.670 -1.730 5.840 -1.560 ;
        RECT 6.030 -1.730 6.200 -1.560 ;
        RECT 6.390 -1.730 6.560 -1.560 ;
        RECT 7.110 -1.730 7.280 -1.560 ;
        RECT 7.470 -1.730 7.640 -1.560 ;
        RECT 7.830 -1.730 8.000 -1.560 ;
        RECT 8.550 -1.730 8.720 -1.560 ;
        RECT 8.930 -1.730 9.100 -1.560 ;
        RECT 8.930 -3.260 9.100 -3.090 ;
        RECT 1.680 -3.690 1.850 -3.520 ;
        RECT 8.930 -4.120 9.100 -3.950 ;
        RECT 1.680 -4.550 1.850 -4.380 ;
        RECT 1.680 -6.590 1.850 -6.420 ;
        RECT 8.930 -7.020 9.100 -6.850 ;
        RECT 1.680 -7.450 1.850 -7.280 ;
        RECT 8.930 -7.880 9.100 -7.710 ;
        RECT 1.680 -9.410 1.850 -9.240 ;
        RECT 2.075 -9.410 2.245 -9.240 ;
        RECT 2.790 -9.410 2.960 -9.240 ;
        RECT 3.150 -9.410 3.320 -9.240 ;
        RECT 3.510 -9.410 3.680 -9.240 ;
        RECT 4.230 -9.410 4.400 -9.240 ;
        RECT 4.590 -9.410 4.760 -9.240 ;
        RECT 4.950 -9.410 5.120 -9.240 ;
        RECT 5.670 -9.410 5.840 -9.240 ;
        RECT 6.030 -9.410 6.200 -9.240 ;
        RECT 6.390 -9.410 6.560 -9.240 ;
        RECT 7.110 -9.410 7.280 -9.240 ;
        RECT 7.470 -9.410 7.640 -9.240 ;
        RECT 7.830 -9.410 8.000 -9.240 ;
        RECT 8.550 -9.410 8.720 -9.240 ;
        RECT 8.930 -9.410 9.100 -9.240 ;
      LAYER met1 ;
        RECT 1.620 -1.760 1.910 -1.530 ;
        RECT 8.870 -1.760 9.160 -1.530 ;
        RECT 1.680 -3.490 1.850 -1.760 ;
        RECT 8.930 -3.060 9.100 -1.760 ;
        RECT 8.900 -3.290 9.130 -3.060 ;
        RECT 1.650 -3.720 1.880 -3.490 ;
        RECT 1.680 -4.350 1.850 -3.720 ;
        RECT 8.930 -3.920 9.100 -3.290 ;
        RECT 8.900 -4.150 9.130 -3.920 ;
        RECT 1.650 -4.580 1.880 -4.350 ;
        RECT 1.680 -6.390 1.850 -4.580 ;
        RECT 1.650 -6.620 1.880 -6.390 ;
        RECT 1.680 -7.250 1.850 -6.620 ;
        RECT 8.930 -6.820 9.100 -4.150 ;
        RECT 8.900 -7.050 9.130 -6.820 ;
        RECT 1.650 -7.480 1.880 -7.250 ;
        RECT 1.680 -9.210 1.850 -7.480 ;
        RECT 8.930 -7.680 9.100 -7.050 ;
        RECT 8.900 -7.910 9.130 -7.680 ;
        RECT 8.930 -9.210 9.100 -7.910 ;
        RECT 1.620 -9.440 1.910 -9.210 ;
        RECT 8.870 -9.440 9.160 -9.210 ;
    END
  END PSUB
  PIN BL[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 -2.240 2.960 -2.070 ;
        RECT 2.790 -8.900 2.960 -8.730 ;
        RECT 2.865 -22.800 3.195 -22.630 ;
      LAYER mcon ;
        RECT 2.945 -22.800 3.115 -22.630 ;
      LAYER met1 ;
        RECT 2.790 -2.040 2.960 -1.905 ;
        RECT 2.730 -2.270 3.020 -2.040 ;
        RECT 2.790 -8.700 2.960 -2.270 ;
        RECT 2.730 -8.930 3.020 -8.700 ;
        RECT 2.790 -10.455 2.960 -8.930 ;
        RECT 2.790 -10.595 3.025 -10.455 ;
        RECT 2.885 -10.895 3.025 -10.595 ;
        RECT 2.885 -11.155 3.205 -10.895 ;
        RECT 2.870 -22.860 3.190 -22.600 ;
      LAYER via ;
        RECT 2.915 -11.155 3.175 -10.895 ;
        RECT 2.900 -22.860 3.160 -22.600 ;
      LAYER met2 ;
        RECT 2.885 -11.155 3.205 -10.895 ;
        RECT 2.985 -22.600 3.125 -11.155 ;
        RECT 2.870 -22.860 3.190 -22.600 ;
    END
  END BL[0]
  PIN BL[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 3.510 -2.240 3.680 -2.070 ;
        RECT 3.510 -8.900 3.680 -8.730 ;
        RECT 3.275 -13.735 3.605 -13.565 ;
      LAYER mcon ;
        RECT 3.355 -13.735 3.525 -13.565 ;
      LAYER met1 ;
        RECT 3.510 -2.040 3.680 -1.905 ;
        RECT 3.450 -2.270 3.740 -2.040 ;
        RECT 3.510 -8.700 3.680 -2.270 ;
        RECT 3.450 -8.930 3.740 -8.700 ;
        RECT 3.510 -10.455 3.680 -8.930 ;
        RECT 3.465 -10.595 3.680 -10.455 ;
        RECT 3.465 -10.895 3.605 -10.595 ;
        RECT 3.345 -11.215 3.605 -10.895 ;
        RECT 3.280 -13.765 3.600 -13.505 ;
      LAYER via ;
        RECT 3.345 -11.185 3.605 -10.925 ;
        RECT 3.310 -13.765 3.570 -13.505 ;
      LAYER met2 ;
        RECT 3.345 -11.215 3.605 -10.895 ;
        RECT 3.345 -13.505 3.485 -11.215 ;
        RECT 3.280 -13.765 3.600 -13.505 ;
    END
  END BL[1]
  PIN BL[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 4.230 -2.240 4.400 -2.070 ;
        RECT 4.230 -8.900 4.400 -8.730 ;
        RECT 4.305 -22.800 4.635 -22.630 ;
      LAYER mcon ;
        RECT 4.385 -22.800 4.555 -22.630 ;
      LAYER met1 ;
        RECT 4.230 -2.040 4.400 -1.905 ;
        RECT 4.170 -2.270 4.460 -2.040 ;
        RECT 4.230 -8.700 4.400 -2.270 ;
        RECT 4.170 -8.930 4.460 -8.700 ;
        RECT 4.230 -10.455 4.400 -8.930 ;
        RECT 4.230 -10.595 4.465 -10.455 ;
        RECT 4.325 -10.895 4.465 -10.595 ;
        RECT 4.325 -11.155 4.645 -10.895 ;
        RECT 4.310 -22.860 4.630 -22.600 ;
      LAYER via ;
        RECT 4.355 -11.155 4.615 -10.895 ;
        RECT 4.340 -22.860 4.600 -22.600 ;
      LAYER met2 ;
        RECT 4.325 -11.155 4.645 -10.895 ;
        RECT 4.425 -22.600 4.565 -11.155 ;
        RECT 4.310 -22.860 4.630 -22.600 ;
    END
  END BL[2]
  PIN BL[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 4.950 -2.240 5.120 -2.070 ;
        RECT 4.950 -8.900 5.120 -8.730 ;
        RECT 4.715 -13.735 5.045 -13.565 ;
      LAYER mcon ;
        RECT 4.795 -13.735 4.965 -13.565 ;
      LAYER met1 ;
        RECT 4.950 -2.040 5.120 -1.905 ;
        RECT 4.890 -2.270 5.180 -2.040 ;
        RECT 4.950 -8.700 5.120 -2.270 ;
        RECT 4.890 -8.930 5.180 -8.700 ;
        RECT 4.950 -10.455 5.120 -8.930 ;
        RECT 4.905 -10.595 5.120 -10.455 ;
        RECT 4.905 -10.895 5.045 -10.595 ;
        RECT 4.785 -11.215 5.045 -10.895 ;
        RECT 4.720 -13.765 5.040 -13.505 ;
      LAYER via ;
        RECT 4.785 -11.185 5.045 -10.925 ;
        RECT 4.750 -13.765 5.010 -13.505 ;
      LAYER met2 ;
        RECT 4.785 -11.215 5.045 -10.895 ;
        RECT 4.785 -13.505 4.925 -11.215 ;
        RECT 4.720 -13.765 5.040 -13.505 ;
    END
  END BL[3]
  PIN BL[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 5.670 -2.240 5.840 -2.070 ;
        RECT 5.670 -8.900 5.840 -8.730 ;
        RECT 5.745 -22.800 6.075 -22.630 ;
      LAYER mcon ;
        RECT 5.825 -22.800 5.995 -22.630 ;
      LAYER met1 ;
        RECT 5.670 -2.040 5.840 -1.905 ;
        RECT 5.610 -2.270 5.900 -2.040 ;
        RECT 5.670 -8.700 5.840 -2.270 ;
        RECT 5.610 -8.930 5.900 -8.700 ;
        RECT 5.670 -10.455 5.840 -8.930 ;
        RECT 5.670 -10.595 5.905 -10.455 ;
        RECT 5.765 -10.895 5.905 -10.595 ;
        RECT 5.765 -11.155 6.085 -10.895 ;
        RECT 5.750 -22.860 6.070 -22.600 ;
      LAYER via ;
        RECT 5.795 -11.155 6.055 -10.895 ;
        RECT 5.780 -22.860 6.040 -22.600 ;
      LAYER met2 ;
        RECT 5.765 -11.155 6.085 -10.895 ;
        RECT 5.865 -22.600 6.005 -11.155 ;
        RECT 5.750 -22.860 6.070 -22.600 ;
    END
  END BL[4]
  PIN BL[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 6.390 -2.240 6.560 -2.070 ;
        RECT 6.390 -8.900 6.560 -8.730 ;
        RECT 6.155 -13.735 6.485 -13.565 ;
      LAYER mcon ;
        RECT 6.235 -13.735 6.405 -13.565 ;
      LAYER met1 ;
        RECT 6.390 -2.040 6.560 -1.905 ;
        RECT 6.330 -2.270 6.620 -2.040 ;
        RECT 6.390 -8.700 6.560 -2.270 ;
        RECT 6.330 -8.930 6.620 -8.700 ;
        RECT 6.390 -10.455 6.560 -8.930 ;
        RECT 6.345 -10.595 6.560 -10.455 ;
        RECT 6.345 -10.895 6.485 -10.595 ;
        RECT 6.225 -11.215 6.485 -10.895 ;
        RECT 6.160 -13.765 6.480 -13.505 ;
      LAYER via ;
        RECT 6.225 -11.185 6.485 -10.925 ;
        RECT 6.190 -13.765 6.450 -13.505 ;
      LAYER met2 ;
        RECT 6.225 -11.215 6.485 -10.895 ;
        RECT 6.225 -13.505 6.365 -11.215 ;
        RECT 6.160 -13.765 6.480 -13.505 ;
    END
  END BL[5]
  PIN BL[6]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 7.110 -2.240 7.280 -2.070 ;
        RECT 7.110 -8.900 7.280 -8.730 ;
        RECT 7.185 -22.800 7.515 -22.630 ;
      LAYER mcon ;
        RECT 7.265 -22.800 7.435 -22.630 ;
      LAYER met1 ;
        RECT 7.110 -2.040 7.280 -1.905 ;
        RECT 7.050 -2.270 7.340 -2.040 ;
        RECT 7.110 -8.700 7.280 -2.270 ;
        RECT 7.050 -8.930 7.340 -8.700 ;
        RECT 7.110 -10.455 7.280 -8.930 ;
        RECT 7.110 -10.595 7.345 -10.455 ;
        RECT 7.205 -10.895 7.345 -10.595 ;
        RECT 7.205 -11.155 7.525 -10.895 ;
        RECT 7.190 -22.860 7.510 -22.600 ;
      LAYER via ;
        RECT 7.235 -11.155 7.495 -10.895 ;
        RECT 7.220 -22.860 7.480 -22.600 ;
      LAYER met2 ;
        RECT 7.205 -11.155 7.525 -10.895 ;
        RECT 7.305 -22.600 7.445 -11.155 ;
        RECT 7.190 -22.860 7.510 -22.600 ;
    END
  END BL[6]
  PIN BL[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 7.830 -2.240 8.000 -2.070 ;
        RECT 7.830 -8.900 8.000 -8.730 ;
        RECT 7.595 -13.735 7.925 -13.565 ;
      LAYER mcon ;
        RECT 7.675 -13.735 7.845 -13.565 ;
      LAYER met1 ;
        RECT 7.830 -2.040 8.000 -1.905 ;
        RECT 7.770 -2.270 8.060 -2.040 ;
        RECT 7.830 -8.700 8.000 -2.270 ;
        RECT 7.770 -8.930 8.060 -8.700 ;
        RECT 7.830 -10.455 8.000 -8.930 ;
        RECT 7.785 -10.595 8.000 -10.455 ;
        RECT 7.785 -10.895 7.925 -10.595 ;
        RECT 7.665 -11.215 7.925 -10.895 ;
        RECT 7.600 -13.765 7.920 -13.505 ;
      LAYER via ;
        RECT 7.665 -11.185 7.925 -10.925 ;
        RECT 7.630 -13.765 7.890 -13.505 ;
      LAYER met2 ;
        RECT 7.665 -11.215 7.925 -10.895 ;
        RECT 7.665 -13.505 7.805 -11.215 ;
        RECT 7.600 -13.765 7.920 -13.505 ;
    END
  END BL[7]
  PIN SSL[0]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -2.625 8.620 -2.455 ;
    END
  END SSL[0]
  PIN WL0[0]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -3.260 2.340 -3.090 ;
    END
  END WL0[0]
  PIN WL0[1]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -3.690 8.620 -3.520 ;
    END
  END WL0[1]
  PIN WL0[2]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -4.120 2.340 -3.950 ;
    END
  END WL0[2]
  PIN WL0[3]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -4.550 8.620 -4.380 ;
    END
  END WL0[3]
  PIN GSL[0]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 2.125 -5.235 2.295 -5.065 ;
    END
  END GSL[0]
  PIN GSL[1]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 2.125 -5.905 2.295 -5.735 ;
    END
  END GSL[1]
  PIN SL
    ANTENNADIFFAREA 1.344000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 -5.570 2.960 -5.400 ;
        RECT 3.510 -5.570 3.680 -5.400 ;
        RECT 4.230 -5.570 4.400 -5.400 ;
        RECT 4.950 -5.570 5.120 -5.400 ;
        RECT 5.670 -5.570 5.840 -5.400 ;
        RECT 6.390 -5.570 6.560 -5.400 ;
        RECT 7.110 -5.570 7.280 -5.400 ;
        RECT 7.830 -5.570 8.000 -5.400 ;
    END
  END SL
  PIN WL1[2]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -7.020 2.340 -6.850 ;
    END
  END WL1[2]
  PIN WL1[3]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -6.590 8.620 -6.420 ;
    END
  END WL1[3]
  PIN WL1[0]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -7.880 2.340 -7.710 ;
    END
  END WL1[0]
  PIN WL1[1]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -7.450 8.620 -7.280 ;
    END
  END WL1[1]
  PIN out_en[0]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.630 -11.140 3.735 -10.970 ;
        RECT 2.630 -11.680 2.800 -11.140 ;
        RECT 2.630 -25.415 3.065 -25.245 ;
      LAYER met1 ;
        RECT 2.585 -11.755 2.845 -11.435 ;
        RECT 2.585 -25.490 2.845 -25.170 ;
      LAYER via ;
        RECT 2.585 -11.725 2.845 -11.465 ;
        RECT 2.585 -25.460 2.845 -25.200 ;
      LAYER met2 ;
        RECT 2.585 -11.755 2.845 -11.435 ;
        RECT 2.585 -25.170 2.725 -11.755 ;
        RECT 2.585 -25.490 2.845 -25.170 ;
    END
  END out_en[0]
  PIN out[1]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 3.270 -11.750 3.440 -11.330 ;
      LAYER mcon ;
        RECT 3.270 -11.625 3.440 -11.455 ;
      LAYER met1 ;
        RECT 3.625 -11.395 3.885 -11.380 ;
        RECT 3.180 -11.685 3.885 -11.395 ;
        RECT 3.625 -11.700 3.885 -11.685 ;
      LAYER via ;
        RECT 3.625 -11.670 3.885 -11.410 ;
      LAYER met2 ;
        RECT 3.625 -11.700 3.885 -11.380 ;
        RECT 3.745 -25.430 3.885 -11.700 ;
    END
  END out[1]
  PIN out[0]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 3.030 -25.055 3.200 -24.635 ;
    END
  END out[0]
  PIN out_en[1]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 4.070 -11.140 5.175 -10.970 ;
        RECT 4.070 -11.680 4.240 -11.140 ;
        RECT 4.070 -25.415 4.505 -25.245 ;
      LAYER met1 ;
        RECT 4.025 -11.755 4.285 -11.435 ;
        RECT 4.025 -25.490 4.285 -25.170 ;
      LAYER via ;
        RECT 4.025 -11.725 4.285 -11.465 ;
        RECT 4.025 -25.460 4.285 -25.200 ;
      LAYER met2 ;
        RECT 4.025 -11.755 4.285 -11.435 ;
        RECT 4.025 -25.170 4.165 -11.755 ;
        RECT 4.025 -25.490 4.285 -25.170 ;
    END
  END out_en[1]
  PIN out[3]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 4.710 -11.750 4.880 -11.330 ;
      LAYER mcon ;
        RECT 4.710 -11.625 4.880 -11.455 ;
      LAYER met1 ;
        RECT 5.065 -11.395 5.325 -11.380 ;
        RECT 4.620 -11.685 5.325 -11.395 ;
        RECT 5.065 -11.700 5.325 -11.685 ;
      LAYER via ;
        RECT 5.065 -11.670 5.325 -11.410 ;
      LAYER met2 ;
        RECT 5.065 -11.700 5.325 -11.380 ;
        RECT 5.185 -25.430 5.325 -11.700 ;
    END
  END out[3]
  PIN out[2]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 4.470 -25.055 4.640 -24.635 ;
    END
  END out[2]
  PIN out_en[2]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 5.510 -11.140 6.615 -10.970 ;
        RECT 5.510 -11.680 5.680 -11.140 ;
        RECT 5.510 -25.415 5.945 -25.245 ;
      LAYER met1 ;
        RECT 5.465 -11.755 5.725 -11.435 ;
        RECT 5.465 -25.490 5.725 -25.170 ;
      LAYER via ;
        RECT 5.465 -11.725 5.725 -11.465 ;
        RECT 5.465 -25.460 5.725 -25.200 ;
      LAYER met2 ;
        RECT 5.465 -11.755 5.725 -11.435 ;
        RECT 5.465 -25.170 5.605 -11.755 ;
        RECT 5.465 -25.490 5.725 -25.170 ;
    END
  END out_en[2]
  PIN out[5]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 6.150 -11.750 6.320 -11.330 ;
      LAYER mcon ;
        RECT 6.150 -11.625 6.320 -11.455 ;
      LAYER met1 ;
        RECT 6.505 -11.395 6.765 -11.380 ;
        RECT 6.060 -11.685 6.765 -11.395 ;
        RECT 6.505 -11.700 6.765 -11.685 ;
      LAYER via ;
        RECT 6.505 -11.670 6.765 -11.410 ;
      LAYER met2 ;
        RECT 6.505 -11.700 6.765 -11.380 ;
        RECT 6.625 -25.430 6.765 -11.700 ;
    END
  END out[5]
  PIN out[4]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 5.910 -25.055 6.080 -24.635 ;
    END
  END out[4]
  PIN out_en[3]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 6.950 -11.140 8.055 -10.970 ;
        RECT 6.950 -11.680 7.120 -11.140 ;
        RECT 6.950 -25.415 7.385 -25.245 ;
      LAYER met1 ;
        RECT 6.905 -11.755 7.165 -11.435 ;
        RECT 6.905 -25.490 7.165 -25.170 ;
      LAYER via ;
        RECT 6.905 -11.725 7.165 -11.465 ;
        RECT 6.905 -25.460 7.165 -25.200 ;
      LAYER met2 ;
        RECT 6.905 -11.755 7.165 -11.435 ;
        RECT 6.905 -25.170 7.045 -11.755 ;
        RECT 6.905 -25.490 7.165 -25.170 ;
    END
  END out_en[3]
  PIN out[7]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 7.590 -11.750 7.760 -11.330 ;
      LAYER mcon ;
        RECT 7.590 -11.625 7.760 -11.455 ;
      LAYER met1 ;
        RECT 7.945 -11.395 8.205 -11.380 ;
        RECT 7.500 -11.685 8.205 -11.395 ;
        RECT 7.945 -11.700 8.205 -11.685 ;
      LAYER via ;
        RECT 7.945 -11.670 8.205 -11.410 ;
      LAYER met2 ;
        RECT 7.945 -11.700 8.205 -11.380 ;
        RECT 8.065 -25.430 8.205 -11.700 ;
    END
  END out[7]
  PIN out[6]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 7.350 -25.055 7.520 -24.635 ;
    END
  END out[6]
  PIN SSL[1]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 8.450 -8.515 8.620 -8.345 ;
    END
  END SSL[1]
  PIN vssd1
    ANTENNADIFFAREA 3.279200 ;
    PORT
      LAYER pwell ;
        RECT 3.100 -11.880 4.085 -11.200 ;
        RECT 4.540 -11.880 5.525 -11.200 ;
        RECT 5.980 -11.880 6.965 -11.200 ;
        RECT 7.420 -11.880 8.405 -11.200 ;
        RECT 3.100 -12.625 3.920 -11.880 ;
        RECT 4.540 -12.625 5.360 -11.880 ;
        RECT 5.980 -12.625 6.800 -11.880 ;
        RECT 7.420 -12.625 8.240 -11.880 ;
        RECT 2.490 -13.305 3.920 -12.625 ;
        RECT 3.930 -13.305 5.360 -12.625 ;
        RECT 5.370 -13.305 6.800 -12.625 ;
        RECT 6.810 -13.305 8.240 -12.625 ;
        RECT 2.765 -15.415 3.705 -13.305 ;
        RECT 4.205 -15.415 5.145 -13.305 ;
        RECT 5.645 -15.415 6.585 -13.305 ;
        RECT 7.085 -15.415 8.025 -13.305 ;
        RECT 2.550 -16.095 3.920 -15.415 ;
        RECT 3.990 -16.095 5.360 -15.415 ;
        RECT 5.430 -16.095 6.800 -15.415 ;
        RECT 6.870 -16.095 8.240 -15.415 ;
        RECT 2.550 -20.950 3.920 -20.270 ;
        RECT 3.990 -20.950 5.360 -20.270 ;
        RECT 5.430 -20.950 6.800 -20.270 ;
        RECT 6.870 -20.950 8.240 -20.270 ;
        RECT 2.765 -23.060 3.705 -20.950 ;
        RECT 4.205 -23.060 5.145 -20.950 ;
        RECT 5.645 -23.060 6.585 -20.950 ;
        RECT 7.085 -23.060 8.025 -20.950 ;
        RECT 2.550 -23.740 3.980 -23.060 ;
        RECT 3.990 -23.740 5.420 -23.060 ;
        RECT 5.430 -23.740 6.860 -23.060 ;
        RECT 6.870 -23.740 8.300 -23.060 ;
        RECT 2.550 -24.505 3.370 -23.740 ;
        RECT 3.990 -24.505 4.810 -23.740 ;
        RECT 5.430 -24.505 6.250 -23.740 ;
        RECT 6.870 -24.505 7.690 -23.740 ;
        RECT 2.385 -25.185 3.370 -24.505 ;
        RECT 3.825 -25.185 4.810 -24.505 ;
        RECT 5.265 -25.185 6.250 -24.505 ;
        RECT 6.705 -25.185 7.690 -24.505 ;
      LAYER li1 ;
        RECT 3.365 -13.965 3.535 -13.905 ;
        RECT 4.805 -13.965 4.975 -13.905 ;
        RECT 6.245 -13.965 6.415 -13.905 ;
        RECT 7.685 -13.965 7.855 -13.905 ;
        RECT 3.345 -14.135 3.535 -13.965 ;
        RECT 4.785 -14.135 4.975 -13.965 ;
        RECT 6.225 -14.135 6.415 -13.965 ;
        RECT 7.665 -14.135 7.855 -13.965 ;
        RECT 3.365 -14.655 3.535 -14.135 ;
        RECT 4.805 -14.655 4.975 -14.135 ;
        RECT 6.245 -14.655 6.415 -14.135 ;
        RECT 7.685 -14.655 7.855 -14.135 ;
        RECT 3.070 -15.275 3.400 -15.105 ;
        RECT 4.510 -15.275 4.840 -15.105 ;
        RECT 5.950 -15.275 6.280 -15.105 ;
        RECT 7.390 -15.275 7.720 -15.105 ;
        RECT 3.150 -15.920 3.320 -15.275 ;
        RECT 4.590 -15.920 4.760 -15.275 ;
        RECT 6.030 -15.920 6.200 -15.275 ;
        RECT 7.470 -15.920 7.640 -15.275 ;
        RECT 3.150 -21.090 3.320 -20.460 ;
        RECT 4.590 -21.090 4.760 -20.460 ;
        RECT 6.030 -21.090 6.200 -20.460 ;
        RECT 7.470 -21.090 7.640 -20.460 ;
        RECT 3.070 -21.260 3.400 -21.090 ;
        RECT 4.510 -21.260 4.840 -21.090 ;
        RECT 5.950 -21.260 6.280 -21.090 ;
        RECT 7.390 -21.260 7.720 -21.090 ;
        RECT 2.935 -22.230 3.105 -21.710 ;
        RECT 4.375 -22.230 4.545 -21.710 ;
        RECT 5.815 -22.230 5.985 -21.710 ;
        RECT 7.255 -22.230 7.425 -21.710 ;
        RECT 2.935 -22.400 3.125 -22.230 ;
        RECT 4.375 -22.400 4.565 -22.230 ;
        RECT 5.815 -22.400 6.005 -22.230 ;
        RECT 7.255 -22.400 7.445 -22.230 ;
        RECT 2.935 -22.460 3.105 -22.400 ;
        RECT 4.375 -22.460 4.545 -22.400 ;
        RECT 5.815 -22.460 5.985 -22.400 ;
        RECT 7.255 -22.460 7.425 -22.400 ;
      LAYER mcon ;
        RECT 3.345 -14.135 3.515 -13.965 ;
        RECT 4.785 -14.135 4.955 -13.965 ;
        RECT 6.225 -14.135 6.395 -13.965 ;
        RECT 7.665 -14.135 7.835 -13.965 ;
        RECT 3.150 -15.275 3.320 -15.105 ;
        RECT 4.590 -15.275 4.760 -15.105 ;
        RECT 6.030 -15.275 6.200 -15.105 ;
        RECT 7.470 -15.275 7.640 -15.105 ;
        RECT 3.150 -21.260 3.320 -21.090 ;
        RECT 4.590 -21.260 4.760 -21.090 ;
        RECT 6.030 -21.260 6.200 -21.090 ;
        RECT 7.470 -21.260 7.640 -21.090 ;
        RECT 2.955 -22.400 3.125 -22.230 ;
        RECT 4.395 -22.400 4.565 -22.230 ;
        RECT 5.835 -22.400 6.005 -22.230 ;
        RECT 7.275 -22.400 7.445 -22.230 ;
      LAYER met1 ;
        RECT 3.315 -14.195 3.545 -13.905 ;
        RECT 4.755 -14.195 4.985 -13.905 ;
        RECT 6.195 -14.195 6.425 -13.905 ;
        RECT 7.635 -14.195 7.865 -13.905 ;
        RECT 3.315 -15.075 3.455 -14.195 ;
        RECT 4.755 -15.075 4.895 -14.195 ;
        RECT 6.195 -15.075 6.335 -14.195 ;
        RECT 7.635 -15.075 7.775 -14.195 ;
        RECT 3.090 -15.120 3.455 -15.075 ;
        RECT 4.530 -15.120 4.895 -15.075 ;
        RECT 5.970 -15.120 6.335 -15.075 ;
        RECT 7.410 -15.120 7.775 -15.075 ;
        RECT 2.515 -15.305 8.555 -15.120 ;
        RECT 8.415 -21.060 8.555 -15.305 ;
        RECT 2.515 -21.245 8.555 -21.060 ;
        RECT 3.015 -21.290 3.380 -21.245 ;
        RECT 4.455 -21.290 4.820 -21.245 ;
        RECT 5.895 -21.290 6.260 -21.245 ;
        RECT 7.335 -21.290 7.700 -21.245 ;
        RECT 3.015 -22.170 3.155 -21.290 ;
        RECT 4.455 -22.170 4.595 -21.290 ;
        RECT 5.895 -22.170 6.035 -21.290 ;
        RECT 7.335 -22.170 7.475 -21.290 ;
        RECT 2.925 -22.460 3.155 -22.170 ;
        RECT 4.365 -22.460 4.595 -22.170 ;
        RECT 5.805 -22.460 6.035 -22.170 ;
        RECT 7.245 -22.460 7.475 -22.170 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 2.860800 ;
    PORT
      LAYER nwell ;
        RECT 2.335 -19.565 8.455 -16.815 ;
      LAYER li1 ;
        RECT 3.150 -18.105 3.320 -17.010 ;
        RECT 4.590 -18.105 4.760 -17.010 ;
        RECT 6.030 -18.105 6.200 -17.010 ;
        RECT 7.470 -18.105 7.640 -17.010 ;
        RECT 2.515 -18.275 8.275 -18.105 ;
        RECT 3.150 -19.370 3.320 -18.275 ;
        RECT 4.590 -19.370 4.760 -18.275 ;
        RECT 6.030 -19.370 6.200 -18.275 ;
        RECT 7.470 -19.370 7.640 -18.275 ;
      LAYER mcon ;
        RECT 3.150 -18.275 3.320 -18.105 ;
        RECT 4.590 -18.275 4.760 -18.105 ;
        RECT 6.030 -18.275 6.200 -18.105 ;
        RECT 7.470 -18.275 7.640 -18.105 ;
      LAYER met1 ;
        RECT 2.515 -18.305 8.275 -18.075 ;
    END
  END vccd1
  PIN sen1
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 3.200 -12.450 3.530 -12.280 ;
        RECT 4.640 -12.450 4.970 -12.280 ;
        RECT 6.080 -12.450 6.410 -12.280 ;
        RECT 7.520 -12.450 7.850 -12.280 ;
        RECT 3.280 -12.465 3.450 -12.450 ;
        RECT 4.720 -12.465 4.890 -12.450 ;
        RECT 6.160 -12.465 6.330 -12.450 ;
        RECT 7.600 -12.465 7.770 -12.450 ;
        RECT 3.020 -23.935 3.190 -23.920 ;
        RECT 4.460 -23.935 4.630 -23.920 ;
        RECT 5.900 -23.935 6.070 -23.920 ;
        RECT 7.340 -23.935 7.510 -23.920 ;
        RECT 2.940 -24.105 3.270 -23.935 ;
        RECT 4.380 -24.105 4.710 -23.935 ;
        RECT 5.820 -24.105 6.150 -23.935 ;
        RECT 7.260 -24.105 7.590 -23.935 ;
      LAYER mcon ;
        RECT 3.020 -24.090 3.190 -23.920 ;
        RECT 4.460 -24.090 4.630 -23.920 ;
        RECT 5.900 -24.090 6.070 -23.920 ;
        RECT 7.340 -24.090 7.510 -23.920 ;
      LAYER met1 ;
        RECT 2.515 -12.495 8.835 -12.265 ;
        RECT 8.695 -23.890 8.835 -12.495 ;
        RECT 2.515 -24.120 8.835 -23.890 ;
    END
  END sen1
  PIN sen2
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 2.800 -11.940 2.970 -11.925 ;
        RECT 4.240 -11.940 4.410 -11.925 ;
        RECT 5.680 -11.940 5.850 -11.925 ;
        RECT 7.120 -11.940 7.290 -11.925 ;
        RECT 2.720 -12.110 3.050 -11.940 ;
        RECT 4.160 -12.110 4.490 -11.940 ;
        RECT 5.600 -12.110 5.930 -11.940 ;
        RECT 7.040 -12.110 7.370 -11.940 ;
        RECT 3.420 -24.445 3.750 -24.275 ;
        RECT 4.860 -24.445 5.190 -24.275 ;
        RECT 6.300 -24.445 6.630 -24.275 ;
        RECT 7.740 -24.445 8.070 -24.275 ;
        RECT 3.500 -24.460 3.670 -24.445 ;
        RECT 4.940 -24.460 5.110 -24.445 ;
        RECT 6.380 -24.460 6.550 -24.445 ;
        RECT 7.820 -24.460 7.990 -24.445 ;
      LAYER mcon ;
        RECT 2.800 -12.095 2.970 -11.925 ;
        RECT 4.240 -12.095 4.410 -11.925 ;
        RECT 5.680 -12.095 5.850 -11.925 ;
        RECT 7.120 -12.095 7.290 -11.925 ;
      LAYER met1 ;
        RECT 2.515 -12.125 9.115 -11.895 ;
        RECT 8.975 -24.260 9.115 -12.125 ;
        RECT 2.515 -24.490 9.115 -24.260 ;
    END
  END sen2
  OBS
      LAYER nwell ;
        RECT 0.000 -1.430 10.790 0.000 ;
        RECT 0.000 -9.540 1.430 -1.430 ;
        RECT 9.360 -9.540 10.790 -1.430 ;
        RECT 0.000 -10.970 10.790 -9.540 ;
      LAYER li1 ;
        RECT 3.160 -0.350 3.330 -0.180 ;
        RECT 4.600 -0.350 4.770 -0.180 ;
        RECT 6.040 -0.350 6.210 -0.180 ;
        RECT 7.480 -0.350 7.650 -0.180 ;
        RECT 3.160 -10.790 3.330 -10.620 ;
        RECT 4.600 -10.790 4.770 -10.620 ;
        RECT 6.040 -10.790 6.210 -10.620 ;
        RECT 7.480 -10.790 7.650 -10.620 ;
        RECT 3.700 -11.455 3.870 -11.330 ;
        RECT 5.140 -11.455 5.310 -11.330 ;
        RECT 6.580 -11.455 6.750 -11.330 ;
        RECT 8.020 -11.455 8.190 -11.330 ;
        RECT 3.670 -11.625 3.870 -11.455 ;
        RECT 5.110 -11.625 5.310 -11.455 ;
        RECT 6.550 -11.625 6.750 -11.455 ;
        RECT 7.990 -11.625 8.190 -11.455 ;
        RECT 3.700 -12.670 3.870 -11.625 ;
        RECT 5.140 -12.670 5.310 -11.625 ;
        RECT 6.580 -12.670 6.750 -11.625 ;
        RECT 8.020 -12.670 8.190 -11.625 ;
        RECT 2.565 -13.050 2.910 -12.880 ;
        RECT 3.150 -13.220 3.320 -12.755 ;
        RECT 3.665 -12.775 3.870 -12.670 ;
        RECT 3.665 -12.800 3.835 -12.775 ;
        RECT 3.580 -13.130 3.835 -12.800 ;
        RECT 4.005 -13.050 4.350 -12.880 ;
        RECT 3.665 -13.175 3.835 -13.130 ;
        RECT 4.590 -13.220 4.760 -12.755 ;
        RECT 5.105 -12.775 5.310 -12.670 ;
        RECT 5.105 -12.800 5.275 -12.775 ;
        RECT 5.020 -13.130 5.275 -12.800 ;
        RECT 5.445 -13.050 5.790 -12.880 ;
        RECT 5.105 -13.175 5.275 -13.130 ;
        RECT 6.030 -13.220 6.200 -12.755 ;
        RECT 6.545 -12.775 6.750 -12.670 ;
        RECT 6.545 -12.800 6.715 -12.775 ;
        RECT 6.460 -13.130 6.715 -12.800 ;
        RECT 6.885 -13.050 7.230 -12.880 ;
        RECT 6.545 -13.175 6.715 -13.130 ;
        RECT 7.470 -13.220 7.640 -12.755 ;
        RECT 7.985 -12.775 8.190 -12.670 ;
        RECT 7.985 -12.800 8.155 -12.775 ;
        RECT 7.900 -13.130 8.155 -12.800 ;
        RECT 7.985 -13.175 8.155 -13.130 ;
        RECT 2.935 -13.390 3.320 -13.220 ;
        RECT 4.375 -13.390 4.760 -13.220 ;
        RECT 5.815 -13.390 6.200 -13.220 ;
        RECT 7.255 -13.390 7.640 -13.220 ;
        RECT 2.935 -14.655 3.105 -13.390 ;
        RECT 4.375 -14.655 4.545 -13.390 ;
        RECT 5.815 -14.655 5.985 -13.390 ;
        RECT 7.255 -14.655 7.425 -13.390 ;
        RECT 2.600 -14.950 2.815 -14.780 ;
        RECT 3.655 -14.950 3.870 -14.780 ;
        RECT 2.600 -15.590 2.770 -14.950 ;
        RECT 3.700 -15.590 3.870 -14.950 ;
        RECT 2.600 -15.920 2.890 -15.590 ;
        RECT 3.580 -15.920 3.870 -15.590 ;
        RECT 2.600 -16.590 2.770 -15.920 ;
        RECT 2.940 -16.170 3.110 -16.090 ;
        RECT 3.700 -16.170 3.870 -15.920 ;
        RECT 2.940 -16.340 3.870 -16.170 ;
        RECT 2.940 -16.420 3.110 -16.340 ;
        RECT 3.360 -16.590 3.530 -16.510 ;
        RECT 2.600 -16.760 3.530 -16.590 ;
        RECT 2.600 -17.060 2.770 -16.760 ;
        RECT 3.360 -16.840 3.530 -16.760 ;
        RECT 2.600 -17.730 2.890 -17.060 ;
        RECT 3.700 -17.140 3.870 -16.340 ;
        RECT 3.500 -17.310 3.870 -17.140 ;
        RECT 3.700 -17.480 3.870 -17.310 ;
        RECT 3.500 -17.650 3.870 -17.480 ;
        RECT 2.600 -17.835 2.770 -17.730 ;
        RECT 3.700 -17.835 3.870 -17.650 ;
        RECT 4.040 -14.950 4.255 -14.780 ;
        RECT 5.095 -14.950 5.310 -14.780 ;
        RECT 4.040 -15.590 4.210 -14.950 ;
        RECT 5.140 -15.590 5.310 -14.950 ;
        RECT 4.040 -15.920 4.330 -15.590 ;
        RECT 5.020 -15.920 5.310 -15.590 ;
        RECT 4.040 -16.590 4.210 -15.920 ;
        RECT 4.380 -16.170 4.550 -16.090 ;
        RECT 5.140 -16.170 5.310 -15.920 ;
        RECT 4.380 -16.340 5.310 -16.170 ;
        RECT 4.380 -16.420 4.550 -16.340 ;
        RECT 4.800 -16.590 4.970 -16.510 ;
        RECT 4.040 -16.760 4.970 -16.590 ;
        RECT 4.040 -17.060 4.210 -16.760 ;
        RECT 4.800 -16.840 4.970 -16.760 ;
        RECT 4.040 -17.730 4.330 -17.060 ;
        RECT 5.140 -17.140 5.310 -16.340 ;
        RECT 4.940 -17.310 5.310 -17.140 ;
        RECT 5.140 -17.480 5.310 -17.310 ;
        RECT 4.940 -17.650 5.310 -17.480 ;
        RECT 4.040 -17.835 4.210 -17.730 ;
        RECT 5.140 -17.835 5.310 -17.650 ;
        RECT 5.480 -14.950 5.695 -14.780 ;
        RECT 6.535 -14.950 6.750 -14.780 ;
        RECT 5.480 -15.590 5.650 -14.950 ;
        RECT 6.580 -15.590 6.750 -14.950 ;
        RECT 5.480 -15.920 5.770 -15.590 ;
        RECT 6.460 -15.920 6.750 -15.590 ;
        RECT 5.480 -16.590 5.650 -15.920 ;
        RECT 5.820 -16.170 5.990 -16.090 ;
        RECT 6.580 -16.170 6.750 -15.920 ;
        RECT 5.820 -16.340 6.750 -16.170 ;
        RECT 5.820 -16.420 5.990 -16.340 ;
        RECT 6.240 -16.590 6.410 -16.510 ;
        RECT 5.480 -16.760 6.410 -16.590 ;
        RECT 5.480 -17.060 5.650 -16.760 ;
        RECT 6.240 -16.840 6.410 -16.760 ;
        RECT 5.480 -17.730 5.770 -17.060 ;
        RECT 6.580 -17.140 6.750 -16.340 ;
        RECT 6.380 -17.310 6.750 -17.140 ;
        RECT 6.580 -17.480 6.750 -17.310 ;
        RECT 6.380 -17.650 6.750 -17.480 ;
        RECT 5.480 -17.835 5.650 -17.730 ;
        RECT 6.580 -17.835 6.750 -17.650 ;
        RECT 6.920 -14.950 7.135 -14.780 ;
        RECT 7.975 -14.950 8.190 -14.780 ;
        RECT 6.920 -15.590 7.090 -14.950 ;
        RECT 8.020 -15.590 8.190 -14.950 ;
        RECT 6.920 -15.920 7.210 -15.590 ;
        RECT 7.900 -15.920 8.190 -15.590 ;
        RECT 6.920 -16.590 7.090 -15.920 ;
        RECT 7.260 -16.170 7.430 -16.090 ;
        RECT 8.020 -16.170 8.190 -15.920 ;
        RECT 7.260 -16.340 8.190 -16.170 ;
        RECT 7.260 -16.420 7.430 -16.340 ;
        RECT 7.680 -16.590 7.850 -16.510 ;
        RECT 6.920 -16.760 7.850 -16.590 ;
        RECT 6.920 -17.060 7.090 -16.760 ;
        RECT 7.680 -16.840 7.850 -16.760 ;
        RECT 6.920 -17.730 7.210 -17.060 ;
        RECT 8.020 -17.140 8.190 -16.340 ;
        RECT 7.820 -17.310 8.190 -17.140 ;
        RECT 8.020 -17.480 8.190 -17.310 ;
        RECT 7.820 -17.650 8.190 -17.480 ;
        RECT 6.920 -17.835 7.090 -17.730 ;
        RECT 8.020 -17.835 8.190 -17.650 ;
        RECT 2.600 -18.730 2.770 -18.545 ;
        RECT 3.700 -18.730 3.870 -18.545 ;
        RECT 2.600 -18.900 2.970 -18.730 ;
        RECT 3.500 -18.900 3.870 -18.730 ;
        RECT 2.600 -19.070 2.770 -18.900 ;
        RECT 3.700 -19.070 3.870 -18.900 ;
        RECT 2.600 -19.240 2.970 -19.070 ;
        RECT 3.500 -19.240 3.870 -19.070 ;
        RECT 2.600 -20.040 2.770 -19.240 ;
        RECT 2.940 -19.620 3.110 -19.540 ;
        RECT 3.700 -19.620 3.870 -19.240 ;
        RECT 2.940 -19.790 3.870 -19.620 ;
        RECT 2.940 -19.870 3.110 -19.790 ;
        RECT 3.360 -20.040 3.530 -19.960 ;
        RECT 2.600 -20.210 3.530 -20.040 ;
        RECT 2.600 -20.525 2.770 -20.210 ;
        RECT 3.360 -20.290 3.530 -20.210 ;
        RECT 3.700 -20.525 3.870 -19.790 ;
        RECT 2.600 -20.695 2.970 -20.525 ;
        RECT 3.500 -20.695 3.870 -20.525 ;
        RECT 2.600 -21.415 2.770 -20.695 ;
        RECT 3.700 -21.415 3.870 -20.695 ;
        RECT 2.600 -21.585 2.815 -21.415 ;
        RECT 3.655 -21.585 3.870 -21.415 ;
        RECT 4.040 -18.730 4.210 -18.545 ;
        RECT 5.140 -18.730 5.310 -18.545 ;
        RECT 4.040 -18.900 4.410 -18.730 ;
        RECT 4.940 -18.900 5.310 -18.730 ;
        RECT 4.040 -19.070 4.210 -18.900 ;
        RECT 5.140 -19.070 5.310 -18.900 ;
        RECT 4.040 -19.240 4.410 -19.070 ;
        RECT 4.940 -19.240 5.310 -19.070 ;
        RECT 4.040 -20.040 4.210 -19.240 ;
        RECT 4.380 -19.620 4.550 -19.540 ;
        RECT 5.140 -19.620 5.310 -19.240 ;
        RECT 4.380 -19.790 5.310 -19.620 ;
        RECT 4.380 -19.870 4.550 -19.790 ;
        RECT 4.800 -20.040 4.970 -19.960 ;
        RECT 4.040 -20.210 4.970 -20.040 ;
        RECT 4.040 -20.525 4.210 -20.210 ;
        RECT 4.800 -20.290 4.970 -20.210 ;
        RECT 5.140 -20.525 5.310 -19.790 ;
        RECT 4.040 -20.695 4.410 -20.525 ;
        RECT 4.940 -20.695 5.310 -20.525 ;
        RECT 4.040 -21.415 4.210 -20.695 ;
        RECT 5.140 -21.415 5.310 -20.695 ;
        RECT 4.040 -21.585 4.255 -21.415 ;
        RECT 5.095 -21.585 5.310 -21.415 ;
        RECT 5.480 -18.730 5.650 -18.545 ;
        RECT 6.580 -18.730 6.750 -18.545 ;
        RECT 5.480 -18.900 5.850 -18.730 ;
        RECT 6.380 -18.900 6.750 -18.730 ;
        RECT 5.480 -19.070 5.650 -18.900 ;
        RECT 6.580 -19.070 6.750 -18.900 ;
        RECT 5.480 -19.240 5.850 -19.070 ;
        RECT 6.380 -19.240 6.750 -19.070 ;
        RECT 5.480 -20.040 5.650 -19.240 ;
        RECT 5.820 -19.620 5.990 -19.540 ;
        RECT 6.580 -19.620 6.750 -19.240 ;
        RECT 5.820 -19.790 6.750 -19.620 ;
        RECT 5.820 -19.870 5.990 -19.790 ;
        RECT 6.240 -20.040 6.410 -19.960 ;
        RECT 5.480 -20.210 6.410 -20.040 ;
        RECT 5.480 -20.525 5.650 -20.210 ;
        RECT 6.240 -20.290 6.410 -20.210 ;
        RECT 6.580 -20.525 6.750 -19.790 ;
        RECT 5.480 -20.695 5.850 -20.525 ;
        RECT 6.380 -20.695 6.750 -20.525 ;
        RECT 5.480 -21.415 5.650 -20.695 ;
        RECT 6.580 -21.415 6.750 -20.695 ;
        RECT 5.480 -21.585 5.695 -21.415 ;
        RECT 6.535 -21.585 6.750 -21.415 ;
        RECT 6.920 -18.730 7.090 -18.545 ;
        RECT 8.020 -18.730 8.190 -18.545 ;
        RECT 6.920 -18.900 7.290 -18.730 ;
        RECT 7.820 -18.900 8.190 -18.730 ;
        RECT 6.920 -19.070 7.090 -18.900 ;
        RECT 8.020 -19.070 8.190 -18.900 ;
        RECT 6.920 -19.240 7.290 -19.070 ;
        RECT 7.820 -19.240 8.190 -19.070 ;
        RECT 6.920 -20.040 7.090 -19.240 ;
        RECT 7.260 -19.620 7.430 -19.540 ;
        RECT 8.020 -19.620 8.190 -19.240 ;
        RECT 7.260 -19.790 8.190 -19.620 ;
        RECT 7.260 -19.870 7.430 -19.790 ;
        RECT 7.680 -20.040 7.850 -19.960 ;
        RECT 6.920 -20.210 7.850 -20.040 ;
        RECT 6.920 -20.525 7.090 -20.210 ;
        RECT 7.680 -20.290 7.850 -20.210 ;
        RECT 8.020 -20.525 8.190 -19.790 ;
        RECT 6.920 -20.695 7.290 -20.525 ;
        RECT 7.820 -20.695 8.190 -20.525 ;
        RECT 6.920 -21.415 7.090 -20.695 ;
        RECT 8.020 -21.415 8.190 -20.695 ;
        RECT 6.920 -21.585 7.135 -21.415 ;
        RECT 7.975 -21.585 8.190 -21.415 ;
        RECT 3.365 -22.975 3.535 -21.710 ;
        RECT 4.805 -22.975 4.975 -21.710 ;
        RECT 6.245 -22.975 6.415 -21.710 ;
        RECT 7.685 -22.975 7.855 -21.710 ;
        RECT 3.150 -23.145 3.535 -22.975 ;
        RECT 4.590 -23.145 4.975 -22.975 ;
        RECT 6.030 -23.145 6.415 -22.975 ;
        RECT 7.470 -23.145 7.855 -22.975 ;
        RECT 2.600 -23.315 2.770 -23.190 ;
        RECT 2.600 -23.485 2.970 -23.315 ;
        RECT 2.600 -25.055 2.770 -23.485 ;
        RECT 3.150 -23.610 3.320 -23.145 ;
        RECT 3.700 -23.315 3.870 -23.190 ;
        RECT 3.560 -23.485 3.870 -23.315 ;
        RECT 3.700 -23.610 3.870 -23.485 ;
        RECT 4.040 -23.315 4.210 -23.190 ;
        RECT 4.040 -23.485 4.410 -23.315 ;
        RECT 4.040 -25.055 4.210 -23.485 ;
        RECT 4.590 -23.610 4.760 -23.145 ;
        RECT 5.140 -23.315 5.310 -23.190 ;
        RECT 5.000 -23.485 5.310 -23.315 ;
        RECT 5.140 -23.610 5.310 -23.485 ;
        RECT 5.480 -23.315 5.650 -23.190 ;
        RECT 5.480 -23.485 5.850 -23.315 ;
        RECT 5.480 -25.055 5.650 -23.485 ;
        RECT 6.030 -23.610 6.200 -23.145 ;
        RECT 6.580 -23.315 6.750 -23.190 ;
        RECT 6.440 -23.485 6.750 -23.315 ;
        RECT 6.580 -23.610 6.750 -23.485 ;
        RECT 6.920 -23.315 7.090 -23.190 ;
        RECT 6.920 -23.485 7.290 -23.315 ;
        RECT 6.920 -25.055 7.090 -23.485 ;
        RECT 7.470 -23.610 7.640 -23.145 ;
        RECT 8.020 -23.315 8.190 -23.190 ;
        RECT 7.880 -23.485 8.190 -23.315 ;
        RECT 8.020 -23.610 8.190 -23.485 ;
      LAYER mcon ;
        RECT 2.615 -13.050 2.785 -12.880 ;
        RECT 3.650 -13.050 3.820 -12.880 ;
        RECT 4.055 -13.050 4.225 -12.880 ;
        RECT 5.090 -13.050 5.260 -12.880 ;
        RECT 5.495 -13.050 5.665 -12.880 ;
        RECT 6.530 -13.050 6.700 -12.880 ;
        RECT 6.935 -13.050 7.105 -12.880 ;
        RECT 7.970 -13.050 8.140 -12.880 ;
        RECT 2.645 -14.950 2.815 -14.780 ;
        RECT 4.085 -14.950 4.255 -14.780 ;
        RECT 5.525 -14.950 5.695 -14.780 ;
        RECT 6.965 -14.950 7.135 -14.780 ;
        RECT 2.645 -21.585 2.815 -21.415 ;
        RECT 4.085 -21.585 4.255 -21.415 ;
        RECT 5.525 -21.585 5.695 -21.415 ;
        RECT 6.965 -21.585 7.135 -21.415 ;
        RECT 2.615 -23.485 2.785 -23.315 ;
        RECT 3.685 -23.485 3.855 -23.315 ;
        RECT 4.055 -23.485 4.225 -23.315 ;
        RECT 5.125 -23.485 5.295 -23.315 ;
        RECT 5.495 -23.485 5.665 -23.315 ;
        RECT 6.565 -23.485 6.735 -23.315 ;
        RECT 6.935 -23.485 7.105 -23.315 ;
        RECT 8.005 -23.485 8.175 -23.315 ;
      LAYER met1 ;
        RECT 2.585 -13.110 2.815 -12.820 ;
        RECT 3.620 -13.110 3.885 -12.820 ;
        RECT 2.585 -14.750 2.725 -13.110 ;
        RECT 3.745 -14.750 3.885 -13.110 ;
        RECT 2.585 -14.980 2.875 -14.750 ;
        RECT 3.595 -14.980 3.885 -14.750 ;
        RECT 4.025 -13.110 4.255 -12.820 ;
        RECT 5.060 -13.110 5.325 -12.820 ;
        RECT 4.025 -14.750 4.165 -13.110 ;
        RECT 5.185 -14.750 5.325 -13.110 ;
        RECT 4.025 -14.980 4.315 -14.750 ;
        RECT 5.035 -14.980 5.325 -14.750 ;
        RECT 5.465 -13.110 5.695 -12.820 ;
        RECT 6.500 -13.110 6.765 -12.820 ;
        RECT 5.465 -14.750 5.605 -13.110 ;
        RECT 6.625 -14.750 6.765 -13.110 ;
        RECT 5.465 -14.980 5.755 -14.750 ;
        RECT 6.475 -14.980 6.765 -14.750 ;
        RECT 6.905 -13.110 7.135 -12.820 ;
        RECT 7.940 -13.110 8.205 -12.820 ;
        RECT 6.905 -14.750 7.045 -13.110 ;
        RECT 8.065 -14.750 8.205 -13.110 ;
        RECT 6.905 -14.980 7.195 -14.750 ;
        RECT 7.915 -14.980 8.205 -14.750 ;
        RECT 2.585 -21.615 2.875 -21.385 ;
        RECT 3.595 -21.615 3.885 -21.385 ;
        RECT 2.585 -23.255 2.725 -21.615 ;
        RECT 3.745 -23.255 3.885 -21.615 ;
        RECT 2.585 -23.545 2.815 -23.255 ;
        RECT 3.655 -23.545 3.885 -23.255 ;
        RECT 4.025 -21.615 4.315 -21.385 ;
        RECT 5.035 -21.615 5.325 -21.385 ;
        RECT 4.025 -23.255 4.165 -21.615 ;
        RECT 5.185 -23.255 5.325 -21.615 ;
        RECT 4.025 -23.545 4.255 -23.255 ;
        RECT 5.095 -23.545 5.325 -23.255 ;
        RECT 5.465 -21.615 5.755 -21.385 ;
        RECT 6.475 -21.615 6.765 -21.385 ;
        RECT 5.465 -23.255 5.605 -21.615 ;
        RECT 6.625 -23.255 6.765 -21.615 ;
        RECT 5.465 -23.545 5.695 -23.255 ;
        RECT 6.535 -23.545 6.765 -23.255 ;
        RECT 6.905 -21.615 7.195 -21.385 ;
        RECT 7.915 -21.615 8.205 -21.385 ;
        RECT 6.905 -23.255 7.045 -21.615 ;
        RECT 8.065 -23.255 8.205 -21.615 ;
        RECT 6.905 -23.545 7.135 -23.255 ;
        RECT 7.975 -23.545 8.205 -23.255 ;
  END
END flash_array_8x8
END LIBRARY

