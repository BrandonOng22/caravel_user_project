VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO flash_array_8x8
  CLASS BLOCK ;
  FOREIGN flash_array_8x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 93.100 BY 500.000 ;
  PIN sen2
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 75.290 -11.940 75.460 -11.925 ;
        RECT 76.730 -11.940 76.900 -11.925 ;
        RECT 78.170 -11.940 78.340 -11.925 ;
        RECT 79.610 -11.940 79.780 -11.925 ;
        RECT 75.210 -12.110 75.540 -11.940 ;
        RECT 76.650 -12.110 76.980 -11.940 ;
        RECT 78.090 -12.110 78.420 -11.940 ;
        RECT 79.530 -12.110 79.860 -11.940 ;
        RECT 75.910 -24.445 76.240 -24.275 ;
        RECT 77.350 -24.445 77.680 -24.275 ;
        RECT 78.790 -24.445 79.120 -24.275 ;
        RECT 80.230 -24.445 80.560 -24.275 ;
        RECT 75.990 -24.460 76.160 -24.445 ;
        RECT 77.430 -24.460 77.600 -24.445 ;
        RECT 78.870 -24.460 79.040 -24.445 ;
        RECT 80.310 -24.460 80.480 -24.445 ;
      LAYER mcon ;
        RECT 75.290 -12.095 75.460 -11.925 ;
        RECT 76.730 -12.095 76.900 -11.925 ;
        RECT 78.170 -12.095 78.340 -11.925 ;
        RECT 79.610 -12.095 79.780 -11.925 ;
      LAYER met1 ;
        RECT 75.005 -12.125 81.605 -11.895 ;
        RECT 81.465 -24.260 81.605 -12.125 ;
        RECT 75.005 -24.490 81.605 -24.260 ;
    END
  END sen2
  PIN sen1
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 75.690 -12.450 76.020 -12.280 ;
        RECT 77.130 -12.450 77.460 -12.280 ;
        RECT 78.570 -12.450 78.900 -12.280 ;
        RECT 80.010 -12.450 80.340 -12.280 ;
        RECT 75.770 -12.465 75.940 -12.450 ;
        RECT 77.210 -12.465 77.380 -12.450 ;
        RECT 78.650 -12.465 78.820 -12.450 ;
        RECT 80.090 -12.465 80.260 -12.450 ;
        RECT 75.510 -23.935 75.680 -23.920 ;
        RECT 76.950 -23.935 77.120 -23.920 ;
        RECT 78.390 -23.935 78.560 -23.920 ;
        RECT 79.830 -23.935 80.000 -23.920 ;
        RECT 75.430 -24.105 75.760 -23.935 ;
        RECT 76.870 -24.105 77.200 -23.935 ;
        RECT 78.310 -24.105 78.640 -23.935 ;
        RECT 79.750 -24.105 80.080 -23.935 ;
      LAYER mcon ;
        RECT 75.510 -24.090 75.680 -23.920 ;
        RECT 76.950 -24.090 77.120 -23.920 ;
        RECT 78.390 -24.090 78.560 -23.920 ;
        RECT 79.830 -24.090 80.000 -23.920 ;
      LAYER met1 ;
        RECT 75.005 -12.495 81.325 -12.265 ;
        RECT 81.185 -23.890 81.325 -12.495 ;
        RECT 75.005 -24.120 81.325 -23.890 ;
    END
  END sen1
  PIN BL[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 80.240 -2.240 80.570 -2.070 ;
        RECT 80.240 -8.900 80.570 -8.730 ;
        RECT 80.085 -13.735 80.415 -13.565 ;
      LAYER mcon ;
        RECT 80.320 -2.240 80.490 -2.070 ;
        RECT 80.320 -8.900 80.490 -8.730 ;
        RECT 80.165 -13.735 80.335 -13.565 ;
      LAYER met1 ;
        RECT 80.320 -2.040 80.490 -1.905 ;
        RECT 80.260 -2.270 80.550 -2.040 ;
        RECT 80.320 -8.700 80.490 -2.270 ;
        RECT 80.260 -8.930 80.550 -8.700 ;
        RECT 80.320 -10.455 80.490 -8.930 ;
        RECT 80.275 -10.595 80.490 -10.455 ;
        RECT 80.275 -10.895 80.415 -10.595 ;
        RECT 80.155 -11.215 80.415 -10.895 ;
        RECT 80.090 -13.765 80.410 -13.505 ;
      LAYER via ;
        RECT 80.155 -11.185 80.415 -10.925 ;
        RECT 80.120 -13.765 80.380 -13.505 ;
      LAYER met2 ;
        RECT 80.155 -11.215 80.415 -10.895 ;
        RECT 80.155 -13.505 80.295 -11.215 ;
        RECT 80.090 -13.765 80.410 -13.505 ;
    END
  END BL[7]
  PIN BL[6]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 79.520 -2.240 79.850 -2.070 ;
        RECT 79.520 -8.900 79.850 -8.730 ;
        RECT 79.675 -22.800 80.005 -22.630 ;
      LAYER mcon ;
        RECT 79.600 -2.240 79.770 -2.070 ;
        RECT 79.600 -8.900 79.770 -8.730 ;
        RECT 79.755 -22.800 79.925 -22.630 ;
      LAYER met1 ;
        RECT 79.600 -2.040 79.770 -1.905 ;
        RECT 79.540 -2.270 79.830 -2.040 ;
        RECT 79.600 -8.700 79.770 -2.270 ;
        RECT 79.540 -8.930 79.830 -8.700 ;
        RECT 79.600 -10.455 79.770 -8.930 ;
        RECT 79.600 -10.595 79.835 -10.455 ;
        RECT 79.695 -10.895 79.835 -10.595 ;
        RECT 79.695 -11.155 80.015 -10.895 ;
        RECT 79.680 -22.860 80.000 -22.600 ;
      LAYER via ;
        RECT 79.725 -11.155 79.985 -10.895 ;
        RECT 79.710 -22.860 79.970 -22.600 ;
      LAYER met2 ;
        RECT 79.695 -11.155 80.015 -10.895 ;
        RECT 79.795 -22.600 79.935 -11.155 ;
        RECT 79.680 -22.860 80.000 -22.600 ;
    END
  END BL[6]
  PIN BL[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 78.800 -2.240 79.130 -2.070 ;
        RECT 78.800 -8.900 79.130 -8.730 ;
        RECT 78.645 -13.735 78.975 -13.565 ;
      LAYER mcon ;
        RECT 78.880 -2.240 79.050 -2.070 ;
        RECT 78.880 -8.900 79.050 -8.730 ;
        RECT 78.725 -13.735 78.895 -13.565 ;
      LAYER met1 ;
        RECT 78.880 -2.040 79.050 -1.905 ;
        RECT 78.820 -2.270 79.110 -2.040 ;
        RECT 78.880 -8.700 79.050 -2.270 ;
        RECT 78.820 -8.930 79.110 -8.700 ;
        RECT 78.880 -10.455 79.050 -8.930 ;
        RECT 78.835 -10.595 79.050 -10.455 ;
        RECT 78.835 -10.895 78.975 -10.595 ;
        RECT 78.715 -11.215 78.975 -10.895 ;
        RECT 78.650 -13.765 78.970 -13.505 ;
      LAYER via ;
        RECT 78.715 -11.185 78.975 -10.925 ;
        RECT 78.680 -13.765 78.940 -13.505 ;
      LAYER met2 ;
        RECT 78.715 -11.215 78.975 -10.895 ;
        RECT 78.715 -13.505 78.855 -11.215 ;
        RECT 78.650 -13.765 78.970 -13.505 ;
    END
  END BL[5]
  PIN BL[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 78.080 -2.240 78.410 -2.070 ;
        RECT 78.080 -8.900 78.410 -8.730 ;
        RECT 78.235 -22.800 78.565 -22.630 ;
      LAYER mcon ;
        RECT 78.160 -2.240 78.330 -2.070 ;
        RECT 78.160 -8.900 78.330 -8.730 ;
        RECT 78.315 -22.800 78.485 -22.630 ;
      LAYER met1 ;
        RECT 78.160 -2.040 78.330 -1.905 ;
        RECT 78.100 -2.270 78.390 -2.040 ;
        RECT 78.160 -8.700 78.330 -2.270 ;
        RECT 78.100 -8.930 78.390 -8.700 ;
        RECT 78.160 -10.455 78.330 -8.930 ;
        RECT 78.160 -10.595 78.395 -10.455 ;
        RECT 78.255 -10.895 78.395 -10.595 ;
        RECT 78.255 -11.155 78.575 -10.895 ;
        RECT 78.240 -22.860 78.560 -22.600 ;
      LAYER via ;
        RECT 78.285 -11.155 78.545 -10.895 ;
        RECT 78.270 -22.860 78.530 -22.600 ;
      LAYER met2 ;
        RECT 78.255 -11.155 78.575 -10.895 ;
        RECT 78.355 -22.600 78.495 -11.155 ;
        RECT 78.240 -22.860 78.560 -22.600 ;
    END
  END BL[4]
  PIN BL[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 77.360 -2.240 77.690 -2.070 ;
        RECT 77.360 -8.900 77.690 -8.730 ;
        RECT 77.205 -13.735 77.535 -13.565 ;
      LAYER mcon ;
        RECT 77.440 -2.240 77.610 -2.070 ;
        RECT 77.440 -8.900 77.610 -8.730 ;
        RECT 77.285 -13.735 77.455 -13.565 ;
      LAYER met1 ;
        RECT 77.440 -2.040 77.610 -1.905 ;
        RECT 77.380 -2.270 77.670 -2.040 ;
        RECT 77.440 -8.700 77.610 -2.270 ;
        RECT 77.380 -8.930 77.670 -8.700 ;
        RECT 77.440 -10.455 77.610 -8.930 ;
        RECT 77.395 -10.595 77.610 -10.455 ;
        RECT 77.395 -10.895 77.535 -10.595 ;
        RECT 77.275 -11.215 77.535 -10.895 ;
        RECT 77.210 -13.765 77.530 -13.505 ;
      LAYER via ;
        RECT 77.275 -11.185 77.535 -10.925 ;
        RECT 77.240 -13.765 77.500 -13.505 ;
      LAYER met2 ;
        RECT 77.275 -11.215 77.535 -10.895 ;
        RECT 77.275 -13.505 77.415 -11.215 ;
        RECT 77.210 -13.765 77.530 -13.505 ;
    END
  END BL[3]
  PIN BL[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 76.640 -2.240 76.970 -2.070 ;
        RECT 76.640 -8.900 76.970 -8.730 ;
        RECT 76.795 -22.800 77.125 -22.630 ;
      LAYER mcon ;
        RECT 76.720 -2.240 76.890 -2.070 ;
        RECT 76.720 -8.900 76.890 -8.730 ;
        RECT 76.875 -22.800 77.045 -22.630 ;
      LAYER met1 ;
        RECT 76.720 -2.040 76.890 -1.905 ;
        RECT 76.660 -2.270 76.950 -2.040 ;
        RECT 76.720 -8.700 76.890 -2.270 ;
        RECT 76.660 -8.930 76.950 -8.700 ;
        RECT 76.720 -10.455 76.890 -8.930 ;
        RECT 76.720 -10.595 76.955 -10.455 ;
        RECT 76.815 -10.895 76.955 -10.595 ;
        RECT 76.815 -11.155 77.135 -10.895 ;
        RECT 76.800 -22.860 77.120 -22.600 ;
      LAYER via ;
        RECT 76.845 -11.155 77.105 -10.895 ;
        RECT 76.830 -22.860 77.090 -22.600 ;
      LAYER met2 ;
        RECT 76.815 -11.155 77.135 -10.895 ;
        RECT 76.915 -22.600 77.055 -11.155 ;
        RECT 76.800 -22.860 77.120 -22.600 ;
    END
  END BL[2]
  PIN BL[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 75.920 -2.240 76.250 -2.070 ;
        RECT 75.920 -8.900 76.250 -8.730 ;
        RECT 75.765 -13.735 76.095 -13.565 ;
      LAYER mcon ;
        RECT 76.000 -2.240 76.170 -2.070 ;
        RECT 76.000 -8.900 76.170 -8.730 ;
        RECT 75.845 -13.735 76.015 -13.565 ;
      LAYER met1 ;
        RECT 76.000 -2.040 76.170 -1.905 ;
        RECT 75.940 -2.270 76.230 -2.040 ;
        RECT 76.000 -8.700 76.170 -2.270 ;
        RECT 75.940 -8.930 76.230 -8.700 ;
        RECT 76.000 -10.455 76.170 -8.930 ;
        RECT 75.955 -10.595 76.170 -10.455 ;
        RECT 75.955 -10.895 76.095 -10.595 ;
        RECT 75.835 -11.215 76.095 -10.895 ;
        RECT 75.770 -13.765 76.090 -13.505 ;
      LAYER via ;
        RECT 75.835 -11.185 76.095 -10.925 ;
        RECT 75.800 -13.765 76.060 -13.505 ;
      LAYER met2 ;
        RECT 75.835 -11.215 76.095 -10.895 ;
        RECT 75.835 -13.505 75.975 -11.215 ;
        RECT 75.770 -13.765 76.090 -13.505 ;
    END
  END BL[1]
  PIN BL[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.273000 ;
    PORT
      LAYER li1 ;
        RECT 75.200 -2.240 75.530 -2.070 ;
        RECT 75.200 -8.900 75.530 -8.730 ;
        RECT 75.355 -22.800 75.685 -22.630 ;
      LAYER mcon ;
        RECT 75.280 -2.240 75.450 -2.070 ;
        RECT 75.280 -8.900 75.450 -8.730 ;
        RECT 75.435 -22.800 75.605 -22.630 ;
      LAYER met1 ;
        RECT 75.280 -2.040 75.450 -1.905 ;
        RECT 75.220 -2.270 75.510 -2.040 ;
        RECT 75.280 -8.700 75.450 -2.270 ;
        RECT 75.220 -8.930 75.510 -8.700 ;
        RECT 75.280 -10.455 75.450 -8.930 ;
        RECT 75.280 -10.595 75.515 -10.455 ;
        RECT 75.375 -10.895 75.515 -10.595 ;
        RECT 75.375 -11.155 75.695 -10.895 ;
        RECT 75.360 -22.860 75.680 -22.600 ;
      LAYER via ;
        RECT 75.405 -11.155 75.665 -10.895 ;
        RECT 75.390 -22.860 75.650 -22.600 ;
      LAYER met2 ;
        RECT 75.375 -11.155 75.695 -10.895 ;
        RECT 75.475 -22.600 75.615 -11.155 ;
        RECT 75.360 -22.860 75.680 -22.600 ;
    END
  END BL[0]
  PIN VBPW
    ANTENNADIFFAREA 8.916200 ;
    PORT
      LAYER li1 ;
        RECT 74.090 -1.730 81.670 -1.560 ;
        RECT 81.340 -3.260 81.670 -3.090 ;
        RECT 74.090 -3.690 74.420 -3.520 ;
        RECT 81.340 -4.120 81.670 -3.950 ;
        RECT 74.090 -4.550 74.420 -4.380 ;
        RECT 74.090 -6.590 74.420 -6.420 ;
        RECT 81.340 -7.020 81.670 -6.850 ;
        RECT 74.090 -7.450 74.420 -7.280 ;
        RECT 81.340 -7.880 81.670 -7.710 ;
        RECT 74.090 -9.410 81.670 -9.240 ;
      LAYER mcon ;
        RECT 74.170 -1.730 74.340 -1.560 ;
        RECT 81.420 -1.730 81.590 -1.560 ;
        RECT 81.420 -3.260 81.590 -3.090 ;
        RECT 74.170 -3.690 74.340 -3.520 ;
        RECT 81.420 -4.120 81.590 -3.950 ;
        RECT 74.170 -4.550 74.340 -4.380 ;
        RECT 74.170 -6.590 74.340 -6.420 ;
        RECT 81.420 -7.020 81.590 -6.850 ;
        RECT 74.170 -7.450 74.340 -7.280 ;
        RECT 81.420 -7.880 81.590 -7.710 ;
        RECT 74.170 -9.410 74.340 -9.240 ;
        RECT 81.420 -9.410 81.590 -9.240 ;
      LAYER met1 ;
        RECT 74.110 -1.760 74.400 -1.530 ;
        RECT 81.360 -1.760 81.650 -1.530 ;
        RECT 74.170 -3.490 74.340 -1.760 ;
        RECT 81.420 -3.060 81.590 -1.760 ;
        RECT 81.390 -3.290 81.620 -3.060 ;
        RECT 74.140 -3.720 74.370 -3.490 ;
        RECT 74.170 -4.350 74.340 -3.720 ;
        RECT 81.420 -3.920 81.590 -3.290 ;
        RECT 81.390 -4.150 81.620 -3.920 ;
        RECT 74.140 -4.580 74.370 -4.350 ;
        RECT 74.170 -6.390 74.340 -4.580 ;
        RECT 74.140 -6.620 74.370 -6.390 ;
        RECT 74.170 -7.250 74.340 -6.620 ;
        RECT 81.420 -6.820 81.590 -4.150 ;
        RECT 81.390 -7.050 81.620 -6.820 ;
        RECT 74.140 -7.480 74.370 -7.250 ;
        RECT 74.170 -9.210 74.340 -7.480 ;
        RECT 81.420 -7.680 81.590 -7.050 ;
        RECT 81.390 -7.910 81.620 -7.680 ;
        RECT 81.420 -9.210 81.590 -7.910 ;
        RECT 74.110 -9.440 74.400 -9.210 ;
        RECT 81.360 -9.440 81.650 -9.210 ;
    END
  END VBPW
  PIN SSL[1]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 80.860 -8.515 81.190 -8.345 ;
    END
  END SSL[1]
  PIN out[6]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 79.840 -25.055 80.010 -24.635 ;
    END
  END out[6]
  PIN out[4]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 78.400 -25.055 78.570 -24.635 ;
    END
  END out[4]
  PIN out[2]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 76.960 -25.055 77.130 -24.635 ;
    END
  END out[2]
  PIN out[0]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 75.520 -25.055 75.690 -24.635 ;
    END
  END out[0]
  PIN WL1[1]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 80.865 -7.450 81.195 -7.280 ;
    END
  END WL1[1]
  PIN WL1[0]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 74.575 -7.880 74.905 -7.710 ;
    END
  END WL1[0]
  PIN WL1[3]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 80.865 -6.590 81.195 -6.420 ;
    END
  END WL1[3]
  PIN WL1[2]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 74.575 -7.020 74.905 -6.850 ;
    END
  END WL1[2]
  PIN SL
    ANTENNADIFFAREA 1.344000 ;
    PORT
      LAYER li1 ;
        RECT 75.005 -5.570 80.765 -5.400 ;
    END
  END SL
  PIN GSL[1]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 74.535 -5.905 74.865 -5.735 ;
    END
  END GSL[1]
  PIN GSL[0]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 74.535 -5.235 74.865 -5.065 ;
    END
  END GSL[0]
  PIN WL0[3]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 80.865 -4.550 81.195 -4.380 ;
    END
  END WL0[3]
  PIN WL0[2]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 74.575 -4.120 74.905 -3.950 ;
    END
  END WL0[2]
  PIN WL0[1]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 80.865 -3.690 81.195 -3.520 ;
    END
  END WL0[1]
  PIN WL0[0]
    ANTENNAGATEAREA 0.792000 ;
    PORT
      LAYER li1 ;
        RECT 74.575 -3.260 74.905 -3.090 ;
    END
  END WL0[0]
  PIN SSL[0]
    ANTENNAGATEAREA 1.680000 ;
    PORT
      LAYER li1 ;
        RECT 80.860 -2.625 81.190 -2.455 ;
    END
  END SSL[0]
  PIN out[7]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 80.080 -11.750 80.250 -11.330 ;
      LAYER mcon ;
        RECT 80.080 -11.625 80.250 -11.455 ;
      LAYER met1 ;
        RECT 80.435 -11.395 80.695 -11.380 ;
        RECT 79.990 -11.685 80.695 -11.395 ;
        RECT 80.435 -11.700 80.695 -11.685 ;
      LAYER via ;
        RECT 80.435 -11.670 80.695 -11.410 ;
      LAYER met2 ;
        RECT 80.435 -11.700 80.695 -11.380 ;
        RECT 80.555 -25.430 80.695 -11.700 ;
    END
  END out[7]
  PIN out_en[3]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 79.440 -11.140 80.545 -10.970 ;
        RECT 79.440 -11.680 79.610 -11.140 ;
        RECT 79.440 -25.415 79.875 -25.245 ;
      LAYER met1 ;
        RECT 79.395 -11.755 79.655 -11.435 ;
        RECT 79.395 -25.490 79.655 -25.170 ;
      LAYER via ;
        RECT 79.395 -11.725 79.655 -11.465 ;
        RECT 79.395 -25.460 79.655 -25.200 ;
      LAYER met2 ;
        RECT 79.395 -11.755 79.655 -11.435 ;
        RECT 79.395 -25.170 79.535 -11.755 ;
        RECT 79.395 -25.490 79.655 -25.170 ;
    END
  END out_en[3]
  PIN out[5]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 78.640 -11.750 78.810 -11.330 ;
      LAYER mcon ;
        RECT 78.640 -11.625 78.810 -11.455 ;
      LAYER met1 ;
        RECT 78.995 -11.395 79.255 -11.380 ;
        RECT 78.550 -11.685 79.255 -11.395 ;
        RECT 78.995 -11.700 79.255 -11.685 ;
      LAYER via ;
        RECT 78.995 -11.670 79.255 -11.410 ;
      LAYER met2 ;
        RECT 78.995 -11.700 79.255 -11.380 ;
        RECT 79.115 -25.430 79.255 -11.700 ;
    END
  END out[5]
  PIN out_en[2]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 78.000 -11.140 79.105 -10.970 ;
        RECT 78.000 -11.680 78.170 -11.140 ;
        RECT 78.000 -25.415 78.435 -25.245 ;
      LAYER met1 ;
        RECT 77.955 -11.755 78.215 -11.435 ;
        RECT 77.955 -25.490 78.215 -25.170 ;
      LAYER via ;
        RECT 77.955 -11.725 78.215 -11.465 ;
        RECT 77.955 -25.460 78.215 -25.200 ;
      LAYER met2 ;
        RECT 77.955 -11.755 78.215 -11.435 ;
        RECT 77.955 -25.170 78.095 -11.755 ;
        RECT 77.955 -25.490 78.215 -25.170 ;
    END
  END out_en[2]
  PIN out[3]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 77.200 -11.750 77.370 -11.330 ;
      LAYER mcon ;
        RECT 77.200 -11.625 77.370 -11.455 ;
      LAYER met1 ;
        RECT 77.555 -11.395 77.815 -11.380 ;
        RECT 77.110 -11.685 77.815 -11.395 ;
        RECT 77.555 -11.700 77.815 -11.685 ;
      LAYER via ;
        RECT 77.555 -11.670 77.815 -11.410 ;
      LAYER met2 ;
        RECT 77.555 -11.700 77.815 -11.380 ;
        RECT 77.675 -25.430 77.815 -11.700 ;
    END
  END out[3]
  PIN out_en[1]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 76.560 -11.140 77.665 -10.970 ;
        RECT 76.560 -11.680 76.730 -11.140 ;
        RECT 76.560 -25.415 76.995 -25.245 ;
      LAYER met1 ;
        RECT 76.515 -11.755 76.775 -11.435 ;
        RECT 76.515 -25.490 76.775 -25.170 ;
      LAYER via ;
        RECT 76.515 -11.725 76.775 -11.465 ;
        RECT 76.515 -25.460 76.775 -25.200 ;
      LAYER met2 ;
        RECT 76.515 -11.755 76.775 -11.435 ;
        RECT 76.515 -25.170 76.655 -11.755 ;
        RECT 76.515 -25.490 76.775 -25.170 ;
    END
  END out_en[1]
  PIN out[1]
    ANTENNADIFFAREA 0.111300 ;
    PORT
      LAYER li1 ;
        RECT 75.760 -11.750 75.930 -11.330 ;
      LAYER mcon ;
        RECT 75.760 -11.625 75.930 -11.455 ;
      LAYER met1 ;
        RECT 76.115 -11.395 76.375 -11.380 ;
        RECT 75.670 -11.685 76.375 -11.395 ;
        RECT 76.115 -11.700 76.375 -11.685 ;
      LAYER via ;
        RECT 76.115 -11.670 76.375 -11.410 ;
      LAYER met2 ;
        RECT 76.115 -11.700 76.375 -11.380 ;
        RECT 76.235 -25.430 76.375 -11.700 ;
    END
  END out[1]
  PIN out_en[0]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 75.120 -11.140 76.225 -10.970 ;
        RECT 75.120 -11.680 75.290 -11.140 ;
        RECT 75.120 -25.415 75.555 -25.245 ;
      LAYER met1 ;
        RECT 75.075 -11.755 75.335 -11.435 ;
        RECT 75.075 -25.490 75.335 -25.170 ;
      LAYER via ;
        RECT 75.075 -11.725 75.335 -11.465 ;
        RECT 75.075 -25.460 75.335 -25.200 ;
      LAYER met2 ;
        RECT 75.075 -11.755 75.335 -11.435 ;
        RECT 75.075 -25.170 75.215 -11.755 ;
        RECT 75.075 -25.490 75.335 -25.170 ;
    END
  END out_en[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 74.825 -19.565 80.945 -16.815 ;
      LAYER li1 ;
        RECT 75.640 -18.105 75.810 -17.010 ;
        RECT 77.080 -18.105 77.250 -17.010 ;
        RECT 78.520 -18.105 78.690 -17.010 ;
        RECT 79.960 -18.105 80.130 -17.010 ;
        RECT 75.005 -18.275 80.765 -18.105 ;
        RECT 75.640 -19.370 75.810 -18.275 ;
        RECT 77.080 -19.370 77.250 -18.275 ;
        RECT 78.520 -19.370 78.690 -18.275 ;
        RECT 79.960 -19.370 80.130 -18.275 ;
      LAYER mcon ;
        RECT 75.640 -18.275 75.810 -18.105 ;
        RECT 77.080 -18.275 77.250 -18.105 ;
        RECT 78.520 -18.275 78.690 -18.105 ;
        RECT 79.960 -18.275 80.130 -18.105 ;
      LAYER met1 ;
        RECT 74.615 -18.075 74.935 -18.060 ;
        RECT 74.615 -18.305 80.765 -18.075 ;
        RECT 74.615 -18.320 74.935 -18.305 ;
      LAYER via ;
        RECT 74.645 -18.320 74.905 -18.060 ;
      LAYER met2 ;
        RECT 38.685 -18.120 41.785 -18.050 ;
        RECT 74.615 -18.120 74.935 -18.060 ;
        RECT 38.685 -18.260 74.935 -18.120 ;
        RECT 38.685 -18.330 41.785 -18.260 ;
        RECT 74.615 -18.320 74.935 -18.260 ;
      LAYER via2 ;
        RECT 39.060 -18.330 39.340 -18.050 ;
        RECT 39.460 -18.330 39.740 -18.050 ;
        RECT 39.860 -18.330 40.140 -18.050 ;
        RECT 40.260 -18.330 40.540 -18.050 ;
        RECT 40.660 -18.330 40.940 -18.050 ;
        RECT 41.060 -18.330 41.340 -18.050 ;
        RECT 41.460 -18.330 41.740 -18.050 ;
      LAYER met3 ;
        RECT 38.685 -18.390 41.785 -17.990 ;
      LAYER via3 ;
        RECT 39.040 -18.350 39.360 -18.030 ;
        RECT 39.440 -18.350 39.760 -18.030 ;
        RECT 39.840 -18.350 40.160 -18.030 ;
        RECT 40.240 -18.350 40.560 -18.030 ;
        RECT 40.640 -18.350 40.960 -18.030 ;
        RECT 41.040 -18.350 41.360 -18.030 ;
        RECT 41.440 -18.350 41.760 -18.030 ;
      LAYER met4 ;
        RECT 38.685 -100.000 41.785 400.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 75.855 -13.965 76.025 -13.905 ;
        RECT 77.295 -13.965 77.465 -13.905 ;
        RECT 78.735 -13.965 78.905 -13.905 ;
        RECT 80.175 -13.965 80.345 -13.905 ;
        RECT 75.835 -14.135 76.025 -13.965 ;
        RECT 77.275 -14.135 77.465 -13.965 ;
        RECT 78.715 -14.135 78.905 -13.965 ;
        RECT 80.155 -14.135 80.345 -13.965 ;
        RECT 75.855 -14.655 76.025 -14.135 ;
        RECT 77.295 -14.655 77.465 -14.135 ;
        RECT 78.735 -14.655 78.905 -14.135 ;
        RECT 80.175 -14.655 80.345 -14.135 ;
        RECT 75.560 -15.275 75.890 -15.105 ;
        RECT 77.000 -15.275 77.330 -15.105 ;
        RECT 78.440 -15.275 78.770 -15.105 ;
        RECT 79.880 -15.275 80.210 -15.105 ;
        RECT 75.640 -15.920 75.810 -15.275 ;
        RECT 77.080 -15.920 77.250 -15.275 ;
        RECT 78.520 -15.920 78.690 -15.275 ;
        RECT 79.960 -15.920 80.130 -15.275 ;
        RECT 75.640 -21.090 75.810 -20.460 ;
        RECT 77.080 -21.090 77.250 -20.460 ;
        RECT 78.520 -21.090 78.690 -20.460 ;
        RECT 79.960 -21.090 80.130 -20.460 ;
        RECT 75.560 -21.260 75.890 -21.090 ;
        RECT 77.000 -21.260 77.330 -21.090 ;
        RECT 78.440 -21.260 78.770 -21.090 ;
        RECT 79.880 -21.260 80.210 -21.090 ;
        RECT 75.425 -22.230 75.595 -21.710 ;
        RECT 76.865 -22.230 77.035 -21.710 ;
        RECT 78.305 -22.230 78.475 -21.710 ;
        RECT 79.745 -22.230 79.915 -21.710 ;
        RECT 75.425 -22.400 75.615 -22.230 ;
        RECT 76.865 -22.400 77.055 -22.230 ;
        RECT 78.305 -22.400 78.495 -22.230 ;
        RECT 79.745 -22.400 79.935 -22.230 ;
        RECT 75.425 -22.460 75.595 -22.400 ;
        RECT 76.865 -22.460 77.035 -22.400 ;
        RECT 78.305 -22.460 78.475 -22.400 ;
        RECT 79.745 -22.460 79.915 -22.400 ;
      LAYER mcon ;
        RECT 75.835 -14.135 76.005 -13.965 ;
        RECT 77.275 -14.135 77.445 -13.965 ;
        RECT 78.715 -14.135 78.885 -13.965 ;
        RECT 80.155 -14.135 80.325 -13.965 ;
        RECT 75.640 -15.275 75.810 -15.105 ;
        RECT 77.080 -15.275 77.250 -15.105 ;
        RECT 78.520 -15.275 78.690 -15.105 ;
        RECT 79.960 -15.275 80.130 -15.105 ;
        RECT 75.640 -21.260 75.810 -21.090 ;
        RECT 77.080 -21.260 77.250 -21.090 ;
        RECT 78.520 -21.260 78.690 -21.090 ;
        RECT 79.960 -21.260 80.130 -21.090 ;
        RECT 75.445 -22.400 75.615 -22.230 ;
        RECT 76.885 -22.400 77.055 -22.230 ;
        RECT 78.325 -22.400 78.495 -22.230 ;
        RECT 79.765 -22.400 79.935 -22.230 ;
      LAYER met1 ;
        RECT 75.805 -14.195 76.035 -13.905 ;
        RECT 77.245 -14.195 77.475 -13.905 ;
        RECT 78.685 -14.195 78.915 -13.905 ;
        RECT 80.125 -14.195 80.355 -13.905 ;
        RECT 75.805 -15.075 75.945 -14.195 ;
        RECT 77.245 -15.075 77.385 -14.195 ;
        RECT 78.685 -15.075 78.825 -14.195 ;
        RECT 80.125 -15.075 80.265 -14.195 ;
        RECT 74.615 -15.120 74.935 -15.085 ;
        RECT 75.580 -15.120 75.945 -15.075 ;
        RECT 77.020 -15.120 77.385 -15.075 ;
        RECT 78.460 -15.120 78.825 -15.075 ;
        RECT 79.900 -15.120 80.265 -15.075 ;
        RECT 74.615 -15.305 81.045 -15.120 ;
        RECT 74.615 -15.345 74.935 -15.305 ;
        RECT 80.905 -21.060 81.045 -15.305 ;
        RECT 75.005 -21.245 81.045 -21.060 ;
        RECT 75.505 -21.290 75.870 -21.245 ;
        RECT 76.945 -21.290 77.310 -21.245 ;
        RECT 78.385 -21.290 78.750 -21.245 ;
        RECT 79.825 -21.290 80.190 -21.245 ;
        RECT 75.505 -22.170 75.645 -21.290 ;
        RECT 76.945 -22.170 77.085 -21.290 ;
        RECT 78.385 -22.170 78.525 -21.290 ;
        RECT 79.825 -22.170 79.965 -21.290 ;
        RECT 75.415 -22.460 75.645 -22.170 ;
        RECT 76.855 -22.460 77.085 -22.170 ;
        RECT 78.295 -22.460 78.525 -22.170 ;
        RECT 79.735 -22.460 79.965 -22.170 ;
      LAYER via ;
        RECT 74.645 -15.345 74.905 -15.085 ;
      LAYER met2 ;
        RECT 74.565 -15.355 74.935 -15.075 ;
      LAYER via2 ;
        RECT 74.610 -15.355 74.890 -15.075 ;
      LAYER met3 ;
        RECT 128.685 -15.050 131.785 -15.015 ;
        RECT 74.585 -15.380 131.785 -15.050 ;
        RECT 128.685 -15.415 131.785 -15.380 ;
      LAYER via3 ;
        RECT 128.690 -15.375 129.010 -15.055 ;
        RECT 129.090 -15.375 129.410 -15.055 ;
        RECT 129.490 -15.375 129.810 -15.055 ;
        RECT 129.890 -15.375 130.210 -15.055 ;
        RECT 130.290 -15.375 130.610 -15.055 ;
        RECT 130.690 -15.375 131.010 -15.055 ;
        RECT 131.090 -15.375 131.410 -15.055 ;
      LAYER met4 ;
        RECT 128.685 -100.000 131.785 400.000 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 72.490 -1.430 83.280 0.000 ;
        RECT 72.490 -9.540 73.920 -1.430 ;
        RECT 81.850 -9.540 83.280 -1.430 ;
        RECT 72.490 -10.970 83.280 -9.540 ;
      LAYER li1 ;
        RECT 75.570 -0.350 75.900 -0.180 ;
        RECT 77.010 -0.350 77.340 -0.180 ;
        RECT 78.450 -0.350 78.780 -0.180 ;
        RECT 79.890 -0.350 80.220 -0.180 ;
        RECT 75.570 -10.790 75.900 -10.620 ;
        RECT 77.010 -10.790 77.340 -10.620 ;
        RECT 78.450 -10.790 78.780 -10.620 ;
        RECT 79.890 -10.790 80.220 -10.620 ;
        RECT 76.190 -11.455 76.360 -11.330 ;
        RECT 77.630 -11.455 77.800 -11.330 ;
        RECT 79.070 -11.455 79.240 -11.330 ;
        RECT 80.510 -11.455 80.680 -11.330 ;
        RECT 76.160 -11.625 76.360 -11.455 ;
        RECT 77.600 -11.625 77.800 -11.455 ;
        RECT 79.040 -11.625 79.240 -11.455 ;
        RECT 80.480 -11.625 80.680 -11.455 ;
        RECT 76.190 -12.670 76.360 -11.625 ;
        RECT 77.630 -12.670 77.800 -11.625 ;
        RECT 79.070 -12.670 79.240 -11.625 ;
        RECT 80.510 -12.670 80.680 -11.625 ;
        RECT 75.055 -13.050 75.400 -12.880 ;
        RECT 75.640 -13.220 75.810 -12.755 ;
        RECT 76.155 -12.775 76.360 -12.670 ;
        RECT 76.155 -12.800 76.325 -12.775 ;
        RECT 76.070 -13.130 76.325 -12.800 ;
        RECT 76.495 -13.050 76.840 -12.880 ;
        RECT 76.155 -13.175 76.325 -13.130 ;
        RECT 77.080 -13.220 77.250 -12.755 ;
        RECT 77.595 -12.775 77.800 -12.670 ;
        RECT 77.595 -12.800 77.765 -12.775 ;
        RECT 77.510 -13.130 77.765 -12.800 ;
        RECT 77.935 -13.050 78.280 -12.880 ;
        RECT 77.595 -13.175 77.765 -13.130 ;
        RECT 78.520 -13.220 78.690 -12.755 ;
        RECT 79.035 -12.775 79.240 -12.670 ;
        RECT 79.035 -12.800 79.205 -12.775 ;
        RECT 78.950 -13.130 79.205 -12.800 ;
        RECT 79.375 -13.050 79.720 -12.880 ;
        RECT 79.035 -13.175 79.205 -13.130 ;
        RECT 79.960 -13.220 80.130 -12.755 ;
        RECT 80.475 -12.775 80.680 -12.670 ;
        RECT 80.475 -12.800 80.645 -12.775 ;
        RECT 80.390 -13.130 80.645 -12.800 ;
        RECT 80.475 -13.175 80.645 -13.130 ;
        RECT 75.425 -13.390 75.810 -13.220 ;
        RECT 76.865 -13.390 77.250 -13.220 ;
        RECT 78.305 -13.390 78.690 -13.220 ;
        RECT 79.745 -13.390 80.130 -13.220 ;
        RECT 75.425 -14.655 75.595 -13.390 ;
        RECT 76.865 -14.655 77.035 -13.390 ;
        RECT 78.305 -14.655 78.475 -13.390 ;
        RECT 79.745 -14.655 79.915 -13.390 ;
        RECT 75.090 -14.950 75.305 -14.780 ;
        RECT 76.145 -14.950 76.360 -14.780 ;
        RECT 75.090 -15.590 75.260 -14.950 ;
        RECT 76.190 -15.590 76.360 -14.950 ;
        RECT 75.090 -15.920 75.380 -15.590 ;
        RECT 76.070 -15.920 76.360 -15.590 ;
        RECT 75.090 -16.590 75.260 -15.920 ;
        RECT 75.430 -16.170 75.600 -16.090 ;
        RECT 76.190 -16.170 76.360 -15.920 ;
        RECT 75.430 -16.340 76.360 -16.170 ;
        RECT 75.430 -16.420 75.600 -16.340 ;
        RECT 75.850 -16.590 76.020 -16.510 ;
        RECT 75.090 -16.760 76.020 -16.590 ;
        RECT 75.090 -17.060 75.260 -16.760 ;
        RECT 75.850 -16.840 76.020 -16.760 ;
        RECT 75.090 -17.730 75.380 -17.060 ;
        RECT 76.190 -17.140 76.360 -16.340 ;
        RECT 75.990 -17.310 76.360 -17.140 ;
        RECT 76.190 -17.480 76.360 -17.310 ;
        RECT 75.990 -17.650 76.360 -17.480 ;
        RECT 75.090 -17.835 75.260 -17.730 ;
        RECT 76.190 -17.835 76.360 -17.650 ;
        RECT 76.530 -14.950 76.745 -14.780 ;
        RECT 77.585 -14.950 77.800 -14.780 ;
        RECT 76.530 -15.590 76.700 -14.950 ;
        RECT 77.630 -15.590 77.800 -14.950 ;
        RECT 76.530 -15.920 76.820 -15.590 ;
        RECT 77.510 -15.920 77.800 -15.590 ;
        RECT 76.530 -16.590 76.700 -15.920 ;
        RECT 76.870 -16.170 77.040 -16.090 ;
        RECT 77.630 -16.170 77.800 -15.920 ;
        RECT 76.870 -16.340 77.800 -16.170 ;
        RECT 76.870 -16.420 77.040 -16.340 ;
        RECT 77.290 -16.590 77.460 -16.510 ;
        RECT 76.530 -16.760 77.460 -16.590 ;
        RECT 76.530 -17.060 76.700 -16.760 ;
        RECT 77.290 -16.840 77.460 -16.760 ;
        RECT 76.530 -17.730 76.820 -17.060 ;
        RECT 77.630 -17.140 77.800 -16.340 ;
        RECT 77.430 -17.310 77.800 -17.140 ;
        RECT 77.630 -17.480 77.800 -17.310 ;
        RECT 77.430 -17.650 77.800 -17.480 ;
        RECT 76.530 -17.835 76.700 -17.730 ;
        RECT 77.630 -17.835 77.800 -17.650 ;
        RECT 77.970 -14.950 78.185 -14.780 ;
        RECT 79.025 -14.950 79.240 -14.780 ;
        RECT 77.970 -15.590 78.140 -14.950 ;
        RECT 79.070 -15.590 79.240 -14.950 ;
        RECT 77.970 -15.920 78.260 -15.590 ;
        RECT 78.950 -15.920 79.240 -15.590 ;
        RECT 77.970 -16.590 78.140 -15.920 ;
        RECT 78.310 -16.170 78.480 -16.090 ;
        RECT 79.070 -16.170 79.240 -15.920 ;
        RECT 78.310 -16.340 79.240 -16.170 ;
        RECT 78.310 -16.420 78.480 -16.340 ;
        RECT 78.730 -16.590 78.900 -16.510 ;
        RECT 77.970 -16.760 78.900 -16.590 ;
        RECT 77.970 -17.060 78.140 -16.760 ;
        RECT 78.730 -16.840 78.900 -16.760 ;
        RECT 77.970 -17.730 78.260 -17.060 ;
        RECT 79.070 -17.140 79.240 -16.340 ;
        RECT 78.870 -17.310 79.240 -17.140 ;
        RECT 79.070 -17.480 79.240 -17.310 ;
        RECT 78.870 -17.650 79.240 -17.480 ;
        RECT 77.970 -17.835 78.140 -17.730 ;
        RECT 79.070 -17.835 79.240 -17.650 ;
        RECT 79.410 -14.950 79.625 -14.780 ;
        RECT 80.465 -14.950 80.680 -14.780 ;
        RECT 79.410 -15.590 79.580 -14.950 ;
        RECT 80.510 -15.590 80.680 -14.950 ;
        RECT 79.410 -15.920 79.700 -15.590 ;
        RECT 80.390 -15.920 80.680 -15.590 ;
        RECT 79.410 -16.590 79.580 -15.920 ;
        RECT 79.750 -16.170 79.920 -16.090 ;
        RECT 80.510 -16.170 80.680 -15.920 ;
        RECT 79.750 -16.340 80.680 -16.170 ;
        RECT 79.750 -16.420 79.920 -16.340 ;
        RECT 80.170 -16.590 80.340 -16.510 ;
        RECT 79.410 -16.760 80.340 -16.590 ;
        RECT 79.410 -17.060 79.580 -16.760 ;
        RECT 80.170 -16.840 80.340 -16.760 ;
        RECT 79.410 -17.730 79.700 -17.060 ;
        RECT 80.510 -17.140 80.680 -16.340 ;
        RECT 80.310 -17.310 80.680 -17.140 ;
        RECT 80.510 -17.480 80.680 -17.310 ;
        RECT 80.310 -17.650 80.680 -17.480 ;
        RECT 79.410 -17.835 79.580 -17.730 ;
        RECT 80.510 -17.835 80.680 -17.650 ;
        RECT 75.090 -18.730 75.260 -18.545 ;
        RECT 76.190 -18.730 76.360 -18.545 ;
        RECT 75.090 -18.900 75.460 -18.730 ;
        RECT 75.990 -18.900 76.360 -18.730 ;
        RECT 75.090 -19.070 75.260 -18.900 ;
        RECT 76.190 -19.070 76.360 -18.900 ;
        RECT 75.090 -19.240 75.460 -19.070 ;
        RECT 75.990 -19.240 76.360 -19.070 ;
        RECT 75.090 -20.040 75.260 -19.240 ;
        RECT 75.430 -19.620 75.600 -19.540 ;
        RECT 76.190 -19.620 76.360 -19.240 ;
        RECT 75.430 -19.790 76.360 -19.620 ;
        RECT 75.430 -19.870 75.600 -19.790 ;
        RECT 75.850 -20.040 76.020 -19.960 ;
        RECT 75.090 -20.210 76.020 -20.040 ;
        RECT 75.090 -20.525 75.260 -20.210 ;
        RECT 75.850 -20.290 76.020 -20.210 ;
        RECT 76.190 -20.525 76.360 -19.790 ;
        RECT 75.090 -20.695 75.460 -20.525 ;
        RECT 75.990 -20.695 76.360 -20.525 ;
        RECT 75.090 -21.415 75.260 -20.695 ;
        RECT 76.190 -21.415 76.360 -20.695 ;
        RECT 75.090 -21.585 75.305 -21.415 ;
        RECT 76.145 -21.585 76.360 -21.415 ;
        RECT 76.530 -18.730 76.700 -18.545 ;
        RECT 77.630 -18.730 77.800 -18.545 ;
        RECT 76.530 -18.900 76.900 -18.730 ;
        RECT 77.430 -18.900 77.800 -18.730 ;
        RECT 76.530 -19.070 76.700 -18.900 ;
        RECT 77.630 -19.070 77.800 -18.900 ;
        RECT 76.530 -19.240 76.900 -19.070 ;
        RECT 77.430 -19.240 77.800 -19.070 ;
        RECT 76.530 -20.040 76.700 -19.240 ;
        RECT 76.870 -19.620 77.040 -19.540 ;
        RECT 77.630 -19.620 77.800 -19.240 ;
        RECT 76.870 -19.790 77.800 -19.620 ;
        RECT 76.870 -19.870 77.040 -19.790 ;
        RECT 77.290 -20.040 77.460 -19.960 ;
        RECT 76.530 -20.210 77.460 -20.040 ;
        RECT 76.530 -20.525 76.700 -20.210 ;
        RECT 77.290 -20.290 77.460 -20.210 ;
        RECT 77.630 -20.525 77.800 -19.790 ;
        RECT 76.530 -20.695 76.900 -20.525 ;
        RECT 77.430 -20.695 77.800 -20.525 ;
        RECT 76.530 -21.415 76.700 -20.695 ;
        RECT 77.630 -21.415 77.800 -20.695 ;
        RECT 76.530 -21.585 76.745 -21.415 ;
        RECT 77.585 -21.585 77.800 -21.415 ;
        RECT 77.970 -18.730 78.140 -18.545 ;
        RECT 79.070 -18.730 79.240 -18.545 ;
        RECT 77.970 -18.900 78.340 -18.730 ;
        RECT 78.870 -18.900 79.240 -18.730 ;
        RECT 77.970 -19.070 78.140 -18.900 ;
        RECT 79.070 -19.070 79.240 -18.900 ;
        RECT 77.970 -19.240 78.340 -19.070 ;
        RECT 78.870 -19.240 79.240 -19.070 ;
        RECT 77.970 -20.040 78.140 -19.240 ;
        RECT 78.310 -19.620 78.480 -19.540 ;
        RECT 79.070 -19.620 79.240 -19.240 ;
        RECT 78.310 -19.790 79.240 -19.620 ;
        RECT 78.310 -19.870 78.480 -19.790 ;
        RECT 78.730 -20.040 78.900 -19.960 ;
        RECT 77.970 -20.210 78.900 -20.040 ;
        RECT 77.970 -20.525 78.140 -20.210 ;
        RECT 78.730 -20.290 78.900 -20.210 ;
        RECT 79.070 -20.525 79.240 -19.790 ;
        RECT 77.970 -20.695 78.340 -20.525 ;
        RECT 78.870 -20.695 79.240 -20.525 ;
        RECT 77.970 -21.415 78.140 -20.695 ;
        RECT 79.070 -21.415 79.240 -20.695 ;
        RECT 77.970 -21.585 78.185 -21.415 ;
        RECT 79.025 -21.585 79.240 -21.415 ;
        RECT 79.410 -18.730 79.580 -18.545 ;
        RECT 80.510 -18.730 80.680 -18.545 ;
        RECT 79.410 -18.900 79.780 -18.730 ;
        RECT 80.310 -18.900 80.680 -18.730 ;
        RECT 79.410 -19.070 79.580 -18.900 ;
        RECT 80.510 -19.070 80.680 -18.900 ;
        RECT 79.410 -19.240 79.780 -19.070 ;
        RECT 80.310 -19.240 80.680 -19.070 ;
        RECT 79.410 -20.040 79.580 -19.240 ;
        RECT 79.750 -19.620 79.920 -19.540 ;
        RECT 80.510 -19.620 80.680 -19.240 ;
        RECT 79.750 -19.790 80.680 -19.620 ;
        RECT 79.750 -19.870 79.920 -19.790 ;
        RECT 80.170 -20.040 80.340 -19.960 ;
        RECT 79.410 -20.210 80.340 -20.040 ;
        RECT 79.410 -20.525 79.580 -20.210 ;
        RECT 80.170 -20.290 80.340 -20.210 ;
        RECT 80.510 -20.525 80.680 -19.790 ;
        RECT 79.410 -20.695 79.780 -20.525 ;
        RECT 80.310 -20.695 80.680 -20.525 ;
        RECT 79.410 -21.415 79.580 -20.695 ;
        RECT 80.510 -21.415 80.680 -20.695 ;
        RECT 79.410 -21.585 79.625 -21.415 ;
        RECT 80.465 -21.585 80.680 -21.415 ;
        RECT 75.855 -22.975 76.025 -21.710 ;
        RECT 77.295 -22.975 77.465 -21.710 ;
        RECT 78.735 -22.975 78.905 -21.710 ;
        RECT 80.175 -22.975 80.345 -21.710 ;
        RECT 75.640 -23.145 76.025 -22.975 ;
        RECT 77.080 -23.145 77.465 -22.975 ;
        RECT 78.520 -23.145 78.905 -22.975 ;
        RECT 79.960 -23.145 80.345 -22.975 ;
        RECT 75.090 -23.315 75.260 -23.190 ;
        RECT 75.090 -23.485 75.460 -23.315 ;
        RECT 75.090 -25.055 75.260 -23.485 ;
        RECT 75.640 -23.610 75.810 -23.145 ;
        RECT 76.190 -23.315 76.360 -23.190 ;
        RECT 76.050 -23.485 76.360 -23.315 ;
        RECT 76.190 -23.610 76.360 -23.485 ;
        RECT 76.530 -23.315 76.700 -23.190 ;
        RECT 76.530 -23.485 76.900 -23.315 ;
        RECT 76.530 -25.055 76.700 -23.485 ;
        RECT 77.080 -23.610 77.250 -23.145 ;
        RECT 77.630 -23.315 77.800 -23.190 ;
        RECT 77.490 -23.485 77.800 -23.315 ;
        RECT 77.630 -23.610 77.800 -23.485 ;
        RECT 77.970 -23.315 78.140 -23.190 ;
        RECT 77.970 -23.485 78.340 -23.315 ;
        RECT 77.970 -25.055 78.140 -23.485 ;
        RECT 78.520 -23.610 78.690 -23.145 ;
        RECT 79.070 -23.315 79.240 -23.190 ;
        RECT 78.930 -23.485 79.240 -23.315 ;
        RECT 79.070 -23.610 79.240 -23.485 ;
        RECT 79.410 -23.315 79.580 -23.190 ;
        RECT 79.410 -23.485 79.780 -23.315 ;
        RECT 79.410 -25.055 79.580 -23.485 ;
        RECT 79.960 -23.610 80.130 -23.145 ;
        RECT 80.510 -23.315 80.680 -23.190 ;
        RECT 80.370 -23.485 80.680 -23.315 ;
        RECT 80.510 -23.610 80.680 -23.485 ;
      LAYER mcon ;
        RECT 75.105 -13.050 75.275 -12.880 ;
        RECT 76.140 -13.050 76.310 -12.880 ;
        RECT 76.545 -13.050 76.715 -12.880 ;
        RECT 77.580 -13.050 77.750 -12.880 ;
        RECT 77.985 -13.050 78.155 -12.880 ;
        RECT 79.020 -13.050 79.190 -12.880 ;
        RECT 79.425 -13.050 79.595 -12.880 ;
        RECT 80.460 -13.050 80.630 -12.880 ;
        RECT 75.135 -14.950 75.305 -14.780 ;
        RECT 76.575 -14.950 76.745 -14.780 ;
        RECT 78.015 -14.950 78.185 -14.780 ;
        RECT 79.455 -14.950 79.625 -14.780 ;
        RECT 75.135 -21.585 75.305 -21.415 ;
        RECT 76.575 -21.585 76.745 -21.415 ;
        RECT 78.015 -21.585 78.185 -21.415 ;
        RECT 79.455 -21.585 79.625 -21.415 ;
        RECT 75.105 -23.485 75.275 -23.315 ;
        RECT 76.175 -23.485 76.345 -23.315 ;
        RECT 76.545 -23.485 76.715 -23.315 ;
        RECT 77.615 -23.485 77.785 -23.315 ;
        RECT 77.985 -23.485 78.155 -23.315 ;
        RECT 79.055 -23.485 79.225 -23.315 ;
        RECT 79.425 -23.485 79.595 -23.315 ;
        RECT 80.495 -23.485 80.665 -23.315 ;
      LAYER met1 ;
        RECT 75.075 -13.110 75.305 -12.820 ;
        RECT 76.110 -13.110 76.375 -12.820 ;
        RECT 75.075 -14.750 75.215 -13.110 ;
        RECT 76.235 -14.750 76.375 -13.110 ;
        RECT 75.075 -14.980 75.365 -14.750 ;
        RECT 76.085 -14.980 76.375 -14.750 ;
        RECT 76.515 -13.110 76.745 -12.820 ;
        RECT 77.550 -13.110 77.815 -12.820 ;
        RECT 76.515 -14.750 76.655 -13.110 ;
        RECT 77.675 -14.750 77.815 -13.110 ;
        RECT 76.515 -14.980 76.805 -14.750 ;
        RECT 77.525 -14.980 77.815 -14.750 ;
        RECT 77.955 -13.110 78.185 -12.820 ;
        RECT 78.990 -13.110 79.255 -12.820 ;
        RECT 77.955 -14.750 78.095 -13.110 ;
        RECT 79.115 -14.750 79.255 -13.110 ;
        RECT 77.955 -14.980 78.245 -14.750 ;
        RECT 78.965 -14.980 79.255 -14.750 ;
        RECT 79.395 -13.110 79.625 -12.820 ;
        RECT 80.430 -13.110 80.695 -12.820 ;
        RECT 79.395 -14.750 79.535 -13.110 ;
        RECT 80.555 -14.750 80.695 -13.110 ;
        RECT 79.395 -14.980 79.685 -14.750 ;
        RECT 80.405 -14.980 80.695 -14.750 ;
        RECT 75.075 -21.615 75.365 -21.385 ;
        RECT 76.085 -21.615 76.375 -21.385 ;
        RECT 75.075 -23.255 75.215 -21.615 ;
        RECT 76.235 -23.255 76.375 -21.615 ;
        RECT 75.075 -23.545 75.305 -23.255 ;
        RECT 76.145 -23.545 76.375 -23.255 ;
        RECT 76.515 -21.615 76.805 -21.385 ;
        RECT 77.525 -21.615 77.815 -21.385 ;
        RECT 76.515 -23.255 76.655 -21.615 ;
        RECT 77.675 -23.255 77.815 -21.615 ;
        RECT 76.515 -23.545 76.745 -23.255 ;
        RECT 77.585 -23.545 77.815 -23.255 ;
        RECT 77.955 -21.615 78.245 -21.385 ;
        RECT 78.965 -21.615 79.255 -21.385 ;
        RECT 77.955 -23.255 78.095 -21.615 ;
        RECT 79.115 -23.255 79.255 -21.615 ;
        RECT 77.955 -23.545 78.185 -23.255 ;
        RECT 79.025 -23.545 79.255 -23.255 ;
        RECT 79.395 -21.615 79.685 -21.385 ;
        RECT 80.405 -21.615 80.695 -21.385 ;
        RECT 79.395 -23.255 79.535 -21.615 ;
        RECT 80.555 -23.255 80.695 -21.615 ;
        RECT 79.395 -23.545 79.625 -23.255 ;
        RECT 80.465 -23.545 80.695 -23.255 ;
  END
END flash_array_8x8
END LIBRARY

