magic
tech sky130A
magscale 1 2
timestamp 1645038762
<< locali >>
rect 260849 439875 260883 440113
rect 260757 439841 260883 439875
rect 260757 439603 260791 439841
rect 260941 439654 260975 439773
rect 260757 439569 261007 439603
rect 260973 439382 261007 439569
rect 262261 439552 262447 439586
rect 262261 439492 262295 439552
rect 262413 439509 262447 439552
rect 262689 439509 262723 440181
rect 262413 439475 262723 439509
rect 262229 439280 262263 439331
rect 260849 439195 260990 439210
rect 260481 439176 260990 439195
rect 260481 439161 260883 439176
rect 260481 436611 260515 439161
rect 260996 438974 261030 439093
rect 262292 439090 262539 439124
rect 260996 438719 261030 438836
rect 260849 438617 260990 438630
rect 260573 438596 260990 438617
rect 260573 438583 260883 438596
rect 260573 435931 260607 438583
rect 261005 438441 261039 438510
rect 261125 438345 261159 438906
rect 262505 438787 262539 439090
rect 262261 438753 262447 438787
rect 262261 438702 262295 438753
rect 262413 438719 262447 438753
rect 262413 438685 262631 438719
rect 262292 438510 262539 438544
rect 260849 438311 261159 438345
rect 260849 438243 260883 438311
rect 260757 438209 260883 438243
rect 262229 438243 262263 438314
rect 260757 438039 260791 438209
rect 260757 438005 260883 438039
rect 260849 436815 260883 438005
rect 260941 435863 260975 437801
rect 262505 435047 262539 438510
rect 261178 434989 261251 435023
rect 261466 434989 261527 435023
rect 261754 434989 261895 435023
rect 262042 434989 262171 435023
rect 261217 432327 261251 434989
rect 261493 432123 261527 434989
rect 261861 431987 261895 434989
rect 262137 432055 262171 434989
rect 262597 434843 262631 438685
<< viali >>
rect 262689 440181 262723 440215
rect 260849 440113 260883 440147
rect 260941 439773 260975 439807
rect 262229 439331 262263 439365
rect 260996 439093 261030 439127
rect 260996 438685 261030 438719
rect 260481 436577 260515 436611
rect 261005 438510 261039 438544
rect 262505 438753 262539 438787
rect 262229 438209 262263 438243
rect 260849 436781 260883 436815
rect 260941 437801 260975 437835
rect 260573 435897 260607 435931
rect 260941 435829 260975 435863
rect 262505 435013 262539 435047
rect 261217 432293 261251 432327
rect 261493 432089 261527 432123
rect 262597 434809 262631 434843
rect 262137 432021 262171 432055
rect 261861 431953 261895 431987
<< metal1 >>
rect 266998 700544 267004 700596
rect 267056 700584 267062 700596
rect 316310 700584 316316 700596
rect 267056 700556 316316 700584
rect 267056 700544 267062 700556
rect 316310 700544 316316 700556
rect 316368 700544 316374 700596
rect 261478 700476 261484 700528
rect 261536 700516 261542 700528
rect 381170 700516 381176 700528
rect 261536 700488 381176 700516
rect 261536 700476 261542 700488
rect 381170 700476 381176 700488
rect 381228 700476 381234 700528
rect 261846 700408 261852 700460
rect 261904 700448 261910 700460
rect 446122 700448 446128 700460
rect 261904 700420 446128 700448
rect 261904 700408 261910 700420
rect 446122 700408 446128 700420
rect 446180 700408 446186 700460
rect 263502 700340 263508 700392
rect 263560 700380 263566 700392
rect 510982 700380 510988 700392
rect 263560 700352 510988 700380
rect 263560 700340 263566 700352
rect 510982 700340 510988 700352
rect 511040 700340 511046 700392
rect 263410 700272 263416 700324
rect 263468 700312 263474 700324
rect 575842 700312 575848 700324
rect 263468 700284 575848 700312
rect 263468 700272 263474 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 56778 700136 56784 700188
rect 56836 700176 56842 700188
rect 57882 700176 57888 700188
rect 56836 700148 57888 700176
rect 56836 700136 56842 700148
rect 57882 700136 57888 700148
rect 57940 700136 57946 700188
rect 186498 700136 186504 700188
rect 186556 700176 186562 700188
rect 187602 700176 187608 700188
rect 186556 700148 187608 700176
rect 186556 700136 186562 700148
rect 187602 700136 187608 700148
rect 187660 700136 187666 700188
rect 251450 700068 251456 700120
rect 251508 700108 251514 700120
rect 252462 700108 252468 700120
rect 251508 700080 252468 700108
rect 251508 700068 251514 700080
rect 252462 700068 252468 700080
rect 252520 700068 252526 700120
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 260834 656888 260840 656940
rect 260892 656928 260898 656940
rect 580166 656928 580172 656940
rect 260892 656900 580172 656928
rect 260892 656888 260898 656900
rect 580166 656888 580172 656900
rect 580224 656888 580230 656940
rect 260926 603100 260932 603152
rect 260984 603140 260990 603152
rect 580166 603140 580172 603152
rect 260984 603112 580172 603140
rect 260984 603100 260990 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 261018 550604 261024 550656
rect 261076 550644 261082 550656
rect 580166 550644 580172 550656
rect 261076 550616 580172 550644
rect 261076 550604 261082 550616
rect 580166 550604 580172 550616
rect 580224 550604 580230 550656
rect 261110 496816 261116 496868
rect 261168 496856 261174 496868
rect 580166 496856 580172 496868
rect 261168 496828 580172 496856
rect 261168 496816 261174 496828
rect 580166 496816 580172 496828
rect 580224 496816 580230 496868
rect 261110 445204 261116 445256
rect 261168 445244 261174 445256
rect 261846 445244 261852 445256
rect 261168 445216 261852 445244
rect 261168 445204 261174 445216
rect 261846 445204 261852 445216
rect 261904 445204 261910 445256
rect 261938 444388 261944 444440
rect 261996 444428 262002 444440
rect 580166 444428 580172 444440
rect 261996 444400 580172 444428
rect 261996 444388 262002 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 262677 440215 262735 440221
rect 262677 440181 262689 440215
rect 262723 440212 262735 440215
rect 263410 440212 263416 440224
rect 262723 440184 263416 440212
rect 262723 440181 262735 440184
rect 262677 440175 262735 440181
rect 263410 440172 263416 440184
rect 263468 440172 263474 440224
rect 260837 440147 260895 440153
rect 260837 440113 260849 440147
rect 260883 440144 260895 440147
rect 266998 440144 267004 440156
rect 260883 440116 267004 440144
rect 260883 440113 260895 440116
rect 260837 440107 260895 440113
rect 266998 440104 267004 440116
rect 267056 440104 267062 440156
rect 260834 439968 260840 440020
rect 260892 440008 260898 440020
rect 260892 439980 262168 440008
rect 260892 439968 260898 439980
rect 260926 439900 260932 439952
rect 260984 439940 260990 439952
rect 260984 439912 261984 439940
rect 260984 439900 260990 439912
rect 260929 439807 260987 439813
rect 260929 439804 260941 439807
rect 253906 439776 260941 439804
rect 3786 439696 3792 439748
rect 3844 439736 3850 439748
rect 253906 439736 253934 439776
rect 260929 439773 260941 439776
rect 260975 439773 260987 439807
rect 260929 439767 260987 439773
rect 261018 439764 261024 439816
rect 261076 439804 261082 439816
rect 261076 439776 261892 439804
rect 261076 439764 261082 439776
rect 3844 439708 253934 439736
rect 3844 439696 3850 439708
rect 261386 439696 261392 439748
rect 261444 439736 261450 439748
rect 261444 439708 261708 439736
rect 261444 439696 261450 439708
rect 261680 439586 261708 439708
rect 261864 439569 261892 439776
rect 261956 439569 261984 439912
rect 262140 439586 262168 439980
rect 262217 439365 262275 439371
rect 262217 439340 262229 439365
rect 262263 439340 262275 439365
rect 262214 439288 262220 439340
rect 262272 439288 262278 439340
rect 261018 439133 261024 439136
rect 260984 439127 261024 439133
rect 260984 439093 260996 439127
rect 260984 439087 261024 439093
rect 261018 439084 261024 439087
rect 261076 439084 261082 439136
rect 262490 438784 262496 438796
rect 262451 438756 262496 438784
rect 262490 438744 262496 438756
rect 262548 438744 262554 438796
rect 261018 438725 261024 438728
rect 260984 438719 261024 438725
rect 260984 438685 260996 438719
rect 260984 438679 261024 438685
rect 261018 438676 261024 438679
rect 261076 438676 261082 438728
rect 260993 438544 261051 438550
rect 260993 438510 261005 438544
rect 261039 438541 261051 438544
rect 261039 438524 261064 438541
rect 260993 438504 261024 438510
rect 261018 438472 261024 438504
rect 261076 438472 261082 438524
rect 262217 438243 262275 438249
rect 262217 438209 262229 438243
rect 262263 438209 262275 438243
rect 262217 438203 262275 438209
rect 262232 438036 262260 438203
rect 263502 438036 263508 438048
rect 262232 438008 263508 438036
rect 263502 437996 263508 438008
rect 263560 437996 263566 438048
rect 260929 437835 260987 437841
rect 260929 437801 260941 437835
rect 260975 437832 260987 437835
rect 261018 437832 261024 437844
rect 260975 437804 261024 437832
rect 260975 437801 260987 437804
rect 260929 437795 260987 437801
rect 261018 437792 261024 437804
rect 261076 437792 261082 437844
rect 3694 436772 3700 436824
rect 3752 436812 3758 436824
rect 260837 436815 260895 436821
rect 260837 436812 260849 436815
rect 3752 436784 260849 436812
rect 3752 436772 3758 436784
rect 260837 436781 260849 436784
rect 260883 436781 260895 436815
rect 260837 436775 260895 436781
rect 252462 436704 252468 436756
rect 252520 436744 252526 436756
rect 252520 436716 260834 436744
rect 252520 436704 252526 436716
rect 260806 436688 260834 436716
rect 122742 436636 122748 436688
rect 122800 436676 122806 436688
rect 122800 436648 260604 436676
rect 260806 436648 260840 436688
rect 122800 436636 122806 436648
rect 187602 436568 187608 436620
rect 187660 436608 187666 436620
rect 260469 436611 260527 436617
rect 260469 436608 260481 436611
rect 187660 436580 260481 436608
rect 187660 436568 187666 436580
rect 260469 436577 260481 436580
rect 260515 436577 260527 436611
rect 260469 436571 260527 436577
rect 260576 436540 260604 436648
rect 260834 436636 260840 436648
rect 260892 436636 260898 436688
rect 260926 436540 260932 436552
rect 260576 436512 260932 436540
rect 260926 436500 260932 436512
rect 260984 436500 260990 436552
rect 3510 435888 3516 435940
rect 3568 435928 3574 435940
rect 260561 435931 260619 435937
rect 260561 435928 260573 435931
rect 3568 435900 260573 435928
rect 3568 435888 3574 435900
rect 260561 435897 260573 435900
rect 260607 435897 260619 435931
rect 260561 435891 260619 435897
rect 57882 435820 57888 435872
rect 57940 435860 57946 435872
rect 260929 435863 260987 435869
rect 260929 435860 260941 435863
rect 57940 435832 260941 435860
rect 57940 435820 57946 435832
rect 260929 435829 260941 435832
rect 260975 435829 260987 435863
rect 260929 435823 260987 435829
rect 262030 435276 262036 435328
rect 262088 435276 262094 435328
rect 262048 435199 262076 435276
rect 262324 435112 262352 435125
rect 264330 435112 264336 435124
rect 262324 435084 264336 435112
rect 264330 435072 264336 435084
rect 264388 435072 264394 435124
rect 3418 435004 3424 435056
rect 3476 435044 3482 435056
rect 262493 435047 262551 435053
rect 262493 435044 262505 435047
rect 3476 435016 262505 435044
rect 3476 435004 3482 435016
rect 262493 435013 262505 435016
rect 262539 435013 262551 435047
rect 262493 435007 262551 435013
rect 261754 434936 261760 434988
rect 261812 434976 261818 434988
rect 261812 434948 261970 434976
rect 261812 434936 261818 434948
rect 3602 434800 3608 434852
rect 3660 434840 3666 434852
rect 262585 434843 262643 434849
rect 262585 434840 262597 434843
rect 3660 434812 262597 434840
rect 3660 434800 3666 434812
rect 262585 434809 262597 434812
rect 262631 434809 262643 434843
rect 262585 434803 262643 434809
rect 261110 434732 261116 434784
rect 261168 434772 261174 434784
rect 261386 434772 261392 434784
rect 261168 434744 261392 434772
rect 261168 434732 261174 434744
rect 261386 434732 261392 434744
rect 261444 434732 261450 434784
rect 262030 434732 262036 434784
rect 262088 434772 262094 434784
rect 264238 434772 264244 434784
rect 262088 434744 264244 434772
rect 262088 434732 262094 434744
rect 264238 434732 264244 434744
rect 264296 434732 264302 434784
rect 260834 432624 260840 432676
rect 260892 432664 260898 432676
rect 261294 432664 261300 432676
rect 260892 432636 261300 432664
rect 260892 432624 260898 432636
rect 261294 432624 261300 432636
rect 261352 432624 261358 432676
rect 261205 432327 261263 432333
rect 261205 432293 261217 432327
rect 261251 432324 261263 432327
rect 262122 432324 262128 432336
rect 261251 432296 262128 432324
rect 261251 432293 261263 432296
rect 261205 432287 261263 432293
rect 262122 432284 262128 432296
rect 262180 432284 262186 432336
rect 261202 432148 261208 432200
rect 261260 432188 261266 432200
rect 261662 432188 261668 432200
rect 261260 432160 261668 432188
rect 261260 432148 261266 432160
rect 261662 432148 261668 432160
rect 261720 432148 261726 432200
rect 261481 432123 261539 432129
rect 261481 432089 261493 432123
rect 261527 432120 261539 432123
rect 262030 432120 262036 432132
rect 261527 432092 262036 432120
rect 261527 432089 261539 432092
rect 261481 432083 261539 432089
rect 262030 432080 262036 432092
rect 262088 432080 262094 432132
rect 261662 432012 261668 432064
rect 261720 432052 261726 432064
rect 262125 432055 262183 432061
rect 262125 432052 262137 432055
rect 261720 432024 262137 432052
rect 261720 432012 261726 432024
rect 262125 432021 262137 432024
rect 262171 432021 262183 432055
rect 262125 432015 262183 432021
rect 261849 431987 261907 431993
rect 261849 431953 261861 431987
rect 261895 431984 261907 431987
rect 261938 431984 261944 431996
rect 261895 431956 261944 431984
rect 261895 431953 261907 431956
rect 261849 431947 261907 431953
rect 261938 431944 261944 431956
rect 261996 431944 262002 431996
rect 261478 431400 261484 431452
rect 261536 431440 261542 431452
rect 261754 431440 261760 431452
rect 261536 431412 261760 431440
rect 261536 431400 261542 431412
rect 261754 431400 261760 431412
rect 261812 431400 261818 431452
rect 261018 431264 261024 431316
rect 261076 431304 261082 431316
rect 261754 431304 261760 431316
rect 261076 431276 261760 431304
rect 261076 431264 261082 431276
rect 261754 431264 261760 431276
rect 261812 431264 261818 431316
rect 261018 431128 261024 431180
rect 261076 431168 261082 431180
rect 262214 431168 262220 431180
rect 261076 431140 262220 431168
rect 261076 431128 261082 431140
rect 262214 431128 262220 431140
rect 262272 431128 262278 431180
rect 261386 391892 261392 391944
rect 261444 391932 261450 391944
rect 580166 391932 580172 391944
rect 261444 391904 580172 391932
rect 261444 391892 261450 391904
rect 580166 391892 580172 391904
rect 580224 391892 580230 391944
rect 261294 339396 261300 339448
rect 261352 339436 261358 339448
rect 579982 339436 579988 339448
rect 261352 339408 579988 339436
rect 261352 339396 261358 339408
rect 579982 339396 579988 339408
rect 580040 339396 580046 339448
rect 261018 313216 261024 313268
rect 261076 313256 261082 313268
rect 580166 313256 580172 313268
rect 261076 313228 580172 313256
rect 261076 313216 261082 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 261754 285608 261760 285660
rect 261812 285648 261818 285660
rect 580166 285648 580172 285660
rect 261812 285620 580172 285648
rect 261812 285608 261818 285620
rect 580166 285608 580172 285620
rect 580224 285608 580230 285660
rect 261662 259360 261668 259412
rect 261720 259400 261726 259412
rect 580166 259400 580172 259412
rect 261720 259372 580172 259400
rect 261720 259360 261726 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 261846 219376 261852 219428
rect 261904 219416 261910 219428
rect 580166 219416 580172 219428
rect 261904 219388 580172 219416
rect 261904 219376 261910 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 261478 206932 261484 206984
rect 261536 206972 261542 206984
rect 579798 206972 579804 206984
rect 261536 206944 579804 206972
rect 261536 206932 261542 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 261938 179324 261944 179376
rect 261996 179364 262002 179376
rect 580166 179364 580172 179376
rect 261996 179336 580172 179364
rect 261996 179324 262002 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 261202 166948 261208 167000
rect 261260 166988 261266 167000
rect 580166 166988 580172 167000
rect 261260 166960 580172 166988
rect 261260 166948 261266 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 261570 139340 261576 139392
rect 261628 139380 261634 139392
rect 580166 139380 580172 139392
rect 261628 139352 580172 139380
rect 261628 139340 261634 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 261110 126896 261116 126948
rect 261168 126936 261174 126948
rect 580166 126936 580172 126948
rect 261168 126908 580172 126936
rect 261168 126896 261174 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 262030 100648 262036 100700
rect 262088 100688 262094 100700
rect 580166 100688 580172 100700
rect 262088 100660 580172 100688
rect 262088 100648 262094 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 260926 86912 260932 86964
rect 260984 86952 260990 86964
rect 580166 86952 580172 86964
rect 260984 86924 580172 86952
rect 260984 86912 260990 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 260834 60664 260840 60716
rect 260892 60704 260898 60716
rect 580166 60704 580172 60716
rect 260892 60676 580172 60704
rect 260892 60664 260898 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 264330 46860 264336 46912
rect 264388 46900 264394 46912
rect 580166 46900 580172 46912
rect 264388 46872 580172 46900
rect 264388 46860 264394 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 262122 20612 262128 20664
rect 262180 20652 262186 20664
rect 579982 20652 579988 20664
rect 262180 20624 579988 20652
rect 262180 20612 262186 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 264238 6808 264244 6860
rect 264296 6848 264302 6860
rect 580166 6848 580172 6860
rect 264296 6820 580172 6848
rect 264296 6808 264302 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
<< via1 >>
rect 267004 700544 267056 700596
rect 316316 700544 316368 700596
rect 261484 700476 261536 700528
rect 381176 700476 381228 700528
rect 261852 700408 261904 700460
rect 446128 700408 446180 700460
rect 263508 700340 263560 700392
rect 510988 700340 511040 700392
rect 263416 700272 263468 700324
rect 575848 700272 575900 700324
rect 56784 700136 56836 700188
rect 57888 700136 57940 700188
rect 186504 700136 186556 700188
rect 187608 700136 187660 700188
rect 251456 700068 251508 700120
rect 252468 700068 252520 700120
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 260840 656888 260892 656940
rect 580172 656888 580224 656940
rect 260932 603100 260984 603152
rect 580172 603100 580224 603152
rect 261024 550604 261076 550656
rect 580172 550604 580224 550656
rect 261116 496816 261168 496868
rect 580172 496816 580224 496868
rect 261116 445204 261168 445256
rect 261852 445204 261904 445256
rect 261944 444388 261996 444440
rect 580172 444388 580224 444440
rect 263416 440172 263468 440224
rect 267004 440104 267056 440156
rect 260840 439968 260892 440020
rect 260932 439900 260984 439952
rect 3792 439696 3844 439748
rect 261024 439764 261076 439816
rect 261392 439696 261444 439748
rect 262220 439331 262229 439340
rect 262229 439331 262263 439340
rect 262263 439331 262272 439340
rect 262220 439288 262272 439331
rect 261024 439127 261076 439136
rect 261024 439093 261030 439127
rect 261030 439093 261076 439127
rect 261024 439084 261076 439093
rect 262496 438787 262548 438796
rect 262496 438753 262505 438787
rect 262505 438753 262539 438787
rect 262539 438753 262548 438787
rect 262496 438744 262548 438753
rect 261024 438719 261076 438728
rect 261024 438685 261030 438719
rect 261030 438685 261076 438719
rect 261024 438676 261076 438685
rect 261024 438510 261039 438524
rect 261039 438510 261076 438524
rect 261024 438472 261076 438510
rect 263508 437996 263560 438048
rect 261024 437792 261076 437844
rect 3700 436772 3752 436824
rect 252468 436704 252520 436756
rect 122748 436636 122800 436688
rect 187608 436568 187660 436620
rect 260840 436636 260892 436688
rect 260932 436500 260984 436552
rect 3516 435888 3568 435940
rect 57888 435820 57940 435872
rect 262036 435276 262088 435328
rect 264336 435072 264388 435124
rect 3424 435004 3476 435056
rect 261760 434936 261812 434988
rect 3608 434800 3660 434852
rect 261116 434732 261168 434784
rect 261392 434732 261444 434784
rect 262036 434732 262088 434784
rect 264244 434732 264296 434784
rect 260840 432624 260892 432676
rect 261300 432624 261352 432676
rect 262128 432284 262180 432336
rect 261208 432148 261260 432200
rect 261668 432148 261720 432200
rect 262036 432080 262088 432132
rect 261668 432012 261720 432064
rect 261944 431944 261996 431996
rect 261484 431400 261536 431452
rect 261760 431400 261812 431452
rect 261024 431264 261076 431316
rect 261760 431264 261812 431316
rect 261024 431128 261076 431180
rect 262220 431128 262272 431180
rect 261392 391892 261444 391944
rect 580172 391892 580224 391944
rect 261300 339396 261352 339448
rect 579988 339396 580040 339448
rect 261024 313216 261076 313268
rect 580172 313216 580224 313268
rect 261760 285608 261812 285660
rect 580172 285608 580224 285660
rect 261668 259360 261720 259412
rect 580172 259360 580224 259412
rect 261852 219376 261904 219428
rect 580172 219376 580224 219428
rect 261484 206932 261536 206984
rect 579804 206932 579856 206984
rect 261944 179324 261996 179376
rect 580172 179324 580224 179376
rect 261208 166948 261260 167000
rect 580172 166948 580224 167000
rect 261576 139340 261628 139392
rect 580172 139340 580224 139392
rect 261116 126896 261168 126948
rect 580172 126896 580224 126948
rect 262036 100648 262088 100700
rect 580172 100648 580224 100700
rect 260932 86912 260984 86964
rect 580172 86912 580224 86964
rect 260840 60664 260892 60716
rect 580172 60664 580224 60716
rect 264336 46860 264388 46912
rect 580172 46860 580224 46912
rect 262128 20612 262180 20664
rect 579988 20612 580040 20664
rect 264244 6808 264296 6860
rect 580172 6808 580224 6860
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 56796 700194 56824 703520
rect 56784 700188 56836 700194
rect 56784 700130 56836 700136
rect 57888 700188 57940 700194
rect 57888 700130 57940 700136
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 435062 3464 697303
rect 3514 645144 3570 645153
rect 3514 645079 3570 645088
rect 3528 435946 3556 645079
rect 3606 593056 3662 593065
rect 3606 592991 3662 593000
rect 3516 435940 3568 435946
rect 3516 435882 3568 435888
rect 3424 435056 3476 435062
rect 3424 434998 3476 435004
rect 3620 434858 3648 592991
rect 3698 540832 3754 540841
rect 3698 540767 3754 540776
rect 3712 436830 3740 540767
rect 3790 488744 3846 488753
rect 3790 488679 3846 488688
rect 3804 439754 3832 488679
rect 3792 439748 3844 439754
rect 3792 439690 3844 439696
rect 3700 436824 3752 436830
rect 3700 436766 3752 436772
rect 57900 435878 57928 700130
rect 121656 699718 121684 703520
rect 186516 700194 186544 703520
rect 186504 700188 186556 700194
rect 186504 700130 186556 700136
rect 187608 700188 187660 700194
rect 187608 700130 187660 700136
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 122760 436694 122788 699654
rect 122748 436688 122800 436694
rect 122748 436630 122800 436636
rect 187620 436626 187648 700130
rect 251468 700126 251496 703520
rect 316328 700602 316356 703520
rect 267004 700596 267056 700602
rect 267004 700538 267056 700544
rect 316316 700596 316368 700602
rect 316316 700538 316368 700544
rect 261484 700528 261536 700534
rect 261484 700470 261536 700476
rect 251456 700120 251508 700126
rect 251456 700062 251508 700068
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 252480 436762 252508 700062
rect 260840 656940 260892 656946
rect 260840 656882 260892 656888
rect 260852 440026 260880 656882
rect 260932 603152 260984 603158
rect 260932 603094 260984 603100
rect 260840 440020 260892 440026
rect 260840 439962 260892 439968
rect 260944 439958 260972 603094
rect 261024 550656 261076 550662
rect 261024 550598 261076 550604
rect 260932 439952 260984 439958
rect 260932 439894 260984 439900
rect 261036 439822 261064 550598
rect 261116 496868 261168 496874
rect 261116 496810 261168 496816
rect 261128 460934 261156 496810
rect 261128 460906 261432 460934
rect 261116 445256 261168 445262
rect 261116 445198 261168 445204
rect 261024 439816 261076 439822
rect 261024 439758 261076 439764
rect 261128 439634 261156 445198
rect 261404 439754 261432 460906
rect 261392 439748 261444 439754
rect 261392 439690 261444 439696
rect 261036 439606 261156 439634
rect 261036 439142 261064 439606
rect 261024 439136 261076 439142
rect 261024 439078 261076 439084
rect 261496 438954 261524 700470
rect 261852 700460 261904 700466
rect 261852 700402 261904 700408
rect 261864 445262 261892 700402
rect 263508 700392 263560 700398
rect 263508 700334 263560 700340
rect 263416 700324 263468 700330
rect 263416 700266 263468 700272
rect 261852 445256 261904 445262
rect 261852 445198 261904 445204
rect 261944 444440 261996 444446
rect 261944 444382 261996 444388
rect 261036 438926 261524 438954
rect 261036 438734 261064 438926
rect 261024 438728 261076 438734
rect 261024 438670 261076 438676
rect 261024 438524 261076 438530
rect 261024 438466 261076 438472
rect 260838 438016 260894 438025
rect 260838 437951 260894 437960
rect 252468 436756 252520 436762
rect 252468 436698 252520 436704
rect 260852 436694 260880 437951
rect 261036 437850 261064 438466
rect 261956 438002 261984 444382
rect 263428 440230 263456 700266
rect 263416 440224 263468 440230
rect 263416 440166 263468 440172
rect 262220 439340 262272 439346
rect 262220 439282 262272 439288
rect 262232 438025 262260 439282
rect 262496 438796 262548 438802
rect 262496 438738 262548 438744
rect 261512 437974 261984 438002
rect 262218 438016 262274 438025
rect 261024 437844 261076 437850
rect 261024 437786 261076 437792
rect 261512 437716 261540 437974
rect 262218 437951 262274 437960
rect 261224 437050 261252 437308
rect 261220 437022 261252 437050
rect 260840 436688 260892 436694
rect 260840 436630 260892 436636
rect 260930 436656 260986 436665
rect 187608 436620 187660 436626
rect 260930 436591 260986 436600
rect 187608 436562 187660 436568
rect 260944 436558 260972 436591
rect 260932 436552 260984 436558
rect 260932 436494 260984 436500
rect 57888 435872 57940 435878
rect 57888 435814 57940 435820
rect 261220 435554 261248 437022
rect 262508 436665 262536 438738
rect 263520 438054 263548 700334
rect 267016 440162 267044 700538
rect 381188 700534 381216 703520
rect 381176 700528 381228 700534
rect 381176 700470 381228 700476
rect 446140 700466 446168 703520
rect 446128 700460 446180 700466
rect 446128 700402 446180 700408
rect 511000 700398 511028 703520
rect 510988 700392 511040 700398
rect 510988 700334 511040 700340
rect 575860 700330 575888 703520
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 580170 657384 580226 657393
rect 580170 657319 580226 657328
rect 580184 656946 580212 657319
rect 580172 656940 580224 656946
rect 580172 656882 580224 656888
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 551168 580226 551177
rect 580170 551103 580226 551112
rect 580184 550662 580212 551103
rect 580172 550656 580224 550662
rect 580172 550598 580224 550604
rect 580170 497992 580226 498001
rect 580170 497927 580226 497936
rect 580184 496874 580212 497927
rect 580172 496868 580224 496874
rect 580172 496810 580224 496816
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 267004 440156 267056 440162
rect 267004 440098 267056 440104
rect 263508 438048 263560 438054
rect 263508 437990 263560 437996
rect 262494 436656 262550 436665
rect 262494 436591 262550 436600
rect 261152 435248 261180 435540
rect 261220 435526 261252 435554
rect 261224 435282 261252 435526
rect 261128 435220 261180 435248
rect 261220 435254 261252 435282
rect 261440 435282 261468 435540
rect 262036 435328 262088 435334
rect 261440 435254 261524 435282
rect 262036 435270 262088 435276
rect 261128 435112 261156 435220
rect 261128 435084 261180 435112
rect 260944 434982 261086 435010
rect 3608 434852 3660 434858
rect 3608 434794 3660 434800
rect 260840 432676 260892 432682
rect 260840 432618 260892 432624
rect 260852 60722 260880 432618
rect 260944 86970 260972 434982
rect 261152 434874 261180 435084
rect 261036 434846 261180 434874
rect 261036 431322 261064 434846
rect 261116 434784 261168 434790
rect 261116 434726 261168 434732
rect 261024 431316 261076 431322
rect 261024 431258 261076 431264
rect 261024 431180 261076 431186
rect 261024 431122 261076 431128
rect 261036 313274 261064 431122
rect 261024 313268 261076 313274
rect 261024 313210 261076 313216
rect 261128 126954 261156 434726
rect 261220 432562 261248 435254
rect 261304 434738 261332 434996
rect 261360 434874 261388 434996
rect 261360 434846 261432 434874
rect 261404 434790 261432 434846
rect 261392 434784 261444 434790
rect 261304 434710 261340 434738
rect 261392 434726 261444 434732
rect 261312 432682 261340 434710
rect 261300 432676 261352 432682
rect 261300 432618 261352 432624
rect 261220 432534 261340 432562
rect 261208 432200 261260 432206
rect 261208 432142 261260 432148
rect 261220 167006 261248 432142
rect 261312 339454 261340 432534
rect 261496 431746 261524 435254
rect 261404 431718 261524 431746
rect 261404 391950 261432 431718
rect 261484 431452 261536 431458
rect 261484 431394 261536 431400
rect 261392 391944 261444 391950
rect 261392 391886 261444 391892
rect 261300 339448 261352 339454
rect 261300 339390 261352 339396
rect 261496 206990 261524 431394
rect 261484 206984 261536 206990
rect 261484 206926 261536 206932
rect 261208 167000 261260 167006
rect 261208 166942 261260 166948
rect 261588 139398 261616 435010
rect 261648 434738 261676 434996
rect 261760 434988 261812 434994
rect 261760 434930 261812 434936
rect 261864 434982 261894 435010
rect 261648 434710 261708 434738
rect 261680 432206 261708 434710
rect 261668 432200 261720 432206
rect 261668 432142 261720 432148
rect 261668 432064 261720 432070
rect 261668 432006 261720 432012
rect 261680 259418 261708 432006
rect 261772 431458 261800 434930
rect 261760 431452 261812 431458
rect 261760 431394 261812 431400
rect 261760 431316 261812 431322
rect 261760 431258 261812 431264
rect 261772 285666 261800 431258
rect 261760 285660 261812 285666
rect 261760 285602 261812 285608
rect 261668 259412 261720 259418
rect 261668 259354 261720 259360
rect 261864 219434 261892 434982
rect 262048 434790 262076 435270
rect 264336 435124 264388 435130
rect 264336 435066 264388 435072
rect 262140 434982 262182 435010
rect 262036 434784 262088 434790
rect 262036 434726 262088 434732
rect 262140 432426 262168 434982
rect 264244 434784 264296 434790
rect 264244 434726 264296 434732
rect 262140 432398 262260 432426
rect 262128 432336 262180 432342
rect 262128 432278 262180 432284
rect 262036 432132 262088 432138
rect 262036 432074 262088 432080
rect 261944 431996 261996 432002
rect 261944 431938 261996 431944
rect 261852 219428 261904 219434
rect 261852 219370 261904 219376
rect 261956 179382 261984 431938
rect 261944 179376 261996 179382
rect 261944 179318 261996 179324
rect 261576 139392 261628 139398
rect 261576 139334 261628 139340
rect 261116 126948 261168 126954
rect 261116 126890 261168 126896
rect 262048 100706 262076 432074
rect 262036 100700 262088 100706
rect 262036 100642 262088 100648
rect 260932 86964 260984 86970
rect 260932 86906 260984 86912
rect 260840 60716 260892 60722
rect 260840 60658 260892 60664
rect 262140 20670 262168 432278
rect 262232 431186 262260 432398
rect 262220 431180 262272 431186
rect 262220 431122 262272 431128
rect 262128 20664 262180 20670
rect 262128 20606 262180 20612
rect 264256 6866 264284 434726
rect 264348 46918 264376 435066
rect 580172 391944 580224 391950
rect 580172 391886 580224 391892
rect 580184 391785 580212 391886
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 579988 339448 580040 339454
rect 579988 339390 580040 339396
rect 580000 338609 580028 339390
rect 579986 338600 580042 338609
rect 579986 338535 580042 338544
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 285660 580224 285666
rect 580172 285602 580224 285608
rect 580184 285433 580212 285602
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 264336 46912 264388 46918
rect 264336 46854 264388 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 264244 6860 264296 6866
rect 264244 6802 264296 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 645088 3570 645144
rect 3606 593000 3662 593056
rect 3698 540776 3754 540832
rect 3790 488688 3846 488744
rect 260838 437960 260894 438016
rect 262218 437960 262274 438016
rect 260930 436600 260986 436656
rect 580170 657328 580226 657384
rect 580170 604152 580226 604208
rect 580170 551112 580226 551168
rect 580170 497936 580226 497992
rect 580170 444760 580226 444816
rect 262494 436600 262550 436656
rect 580170 391720 580226 391776
rect 579986 338544 580042 338600
rect 580170 312024 580226 312080
rect 580170 285368 580226 285424
rect 580170 258848 580226 258904
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 580165 657386 580231 657389
rect 583520 657386 584960 657476
rect 580165 657384 584960 657386
rect 580165 657328 580170 657384
rect 580226 657328 584960 657384
rect 580165 657326 584960 657328
rect 580165 657323 580231 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 3509 645146 3575 645149
rect -960 645144 3575 645146
rect -960 645088 3514 645144
rect 3570 645088 3575 645144
rect -960 645086 3575 645088
rect -960 644996 480 645086
rect 3509 645083 3575 645086
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3601 593058 3667 593061
rect -960 593056 3667 593058
rect -960 593000 3606 593056
rect 3662 593000 3667 593056
rect -960 592998 3667 593000
rect -960 592908 480 592998
rect 3601 592995 3667 592998
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 580165 551170 580231 551173
rect 583520 551170 584960 551260
rect 580165 551168 584960 551170
rect 580165 551112 580170 551168
rect 580226 551112 584960 551168
rect 580165 551110 584960 551112
rect 580165 551107 580231 551110
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3693 540834 3759 540837
rect -960 540832 3759 540834
rect -960 540776 3698 540832
rect 3754 540776 3759 540832
rect -960 540774 3759 540776
rect -960 540684 480 540774
rect 3693 540771 3759 540774
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 580165 497994 580231 497997
rect 583520 497994 584960 498084
rect 580165 497992 584960 497994
rect 580165 497936 580170 497992
rect 580226 497936 584960 497992
rect 580165 497934 584960 497936
rect 580165 497931 580231 497934
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect 3785 488746 3851 488749
rect -960 488744 3851 488746
rect -960 488688 3790 488744
rect 3846 488688 3851 488744
rect -960 488686 3851 488688
rect -960 488596 480 488686
rect 3785 488683 3851 488686
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 260833 438018 260899 438021
rect 262213 438018 262279 438021
rect 260833 438016 262279 438018
rect 260833 437960 260838 438016
rect 260894 437960 262218 438016
rect 262274 437960 262279 438016
rect 260833 437958 262279 437960
rect 260833 437955 260899 437958
rect 262213 437955 262279 437958
rect -960 436508 480 436748
rect 260925 436658 260991 436661
rect 262489 436658 262555 436661
rect 260925 436656 262555 436658
rect 260925 436600 260930 436656
rect 260986 436600 262494 436656
rect 262550 436600 262555 436656
rect 260925 436598 262555 436600
rect 260925 436595 260991 436598
rect 262489 436595 262555 436598
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 579981 338602 580047 338605
rect 583520 338602 584960 338692
rect 579981 338600 584960 338602
rect 579981 338544 579986 338600
rect 580042 338544 584960 338600
rect 579981 338542 584960 338544
rect 579981 338539 580047 338542
rect 583520 338452 584960 338542
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214828 480 215068
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136628 480 136868
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6340 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 583520 6476 584960 6566
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use flash_array_8x8  u_flash_array_8x8
timestamp 1645038762
transform 1 0 246057 0 1 440000
box 7737 -20000 26357 80000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
